// 10b inputs to PCA algorithm


// row 0 pixels 0-31 
assign pca_data_in_10b[0][0] = 10'b0;
assign pca_data_in_10b[0][1] = 10'b0;
assign pca_data_in_10b[0][2] = 10'b0;
assign pca_data_in_10b[0][3] = 10'b0;
assign pca_data_in_10b[0][4] = 10'b0;
assign pca_data_in_10b[0][5] = 10'b0;
assign pca_data_in_10b[0][6] = 10'b0;
assign pca_data_in_10b[0][7] = 10'b0;
assign pca_data_in_10b[0][8] = 10'b0;
assign pca_data_in_10b[0][9] = 10'b0;
assign pca_data_in_10b[0][10] = 10'b0;
assign pca_data_in_10b[0][11] = 10'b0;
assign pca_data_in_10b[0][12] = 10'b0;
assign pca_data_in_10b[0][13] = 10'b0;
assign pca_data_in_10b[0][14] = 10'b0;
assign pca_data_in_10b[0][15] = 10'b0;
assign pca_data_in_10b[0][16] = 10'b0;
assign pca_data_in_10b[0][17] = 10'b0;
assign pca_data_in_10b[0][18] = 10'b0;
assign pca_data_in_10b[0][19] = 10'b0;
assign pca_data_in_10b[0][20] = 10'b0;
assign pca_data_in_10b[0][21] = 10'b0;
assign pca_data_in_10b[0][22] = 10'b0;
assign pca_data_in_10b[0][23] = 10'b0;
assign pca_data_in_10b[0][24] = 10'b0;
assign pca_data_in_10b[0][25] = 10'b0;
assign pca_data_in_10b[0][26] = 10'b0;
assign pca_data_in_10b[0][27] = 10'b0;
assign pca_data_in_10b[0][28] = 10'b0;
assign pca_data_in_10b[0][29] = 10'b0;
assign pca_data_in_10b[0][30] = 10'b0;
assign pca_data_in_10b[0][31] = 10'b0;

// row 1 pixels 0-31 
assign pca_data_in_10b[1][0] = 10'b0;
assign pca_data_in_10b[1][1] = 10'b0;
assign pca_data_in_10b[1][2] = 10'b0;
assign pca_data_in_10b[1][3] = 10'b0;
assign pca_data_in_10b[1][4] = 10'b0;
assign pca_data_in_10b[1][5] = 10'b0;
assign pca_data_in_10b[1][6] = 10'b0;
assign pca_data_in_10b[1][7] = 10'b0;
assign pca_data_in_10b[1][8] = 10'b0;
assign pca_data_in_10b[1][9] = 10'b0;
assign pca_data_in_10b[1][10] = 10'b0;
assign pca_data_in_10b[1][11] = 10'b0;
assign pca_data_in_10b[1][12] = 10'b0;
assign pca_data_in_10b[1][13] = 10'b0;
assign pca_data_in_10b[1][14] = 10'b0;
assign pca_data_in_10b[1][15] = 10'b0;
assign pca_data_in_10b[1][16] = 10'b0;
assign pca_data_in_10b[1][17] = 10'b0;
assign pca_data_in_10b[1][18] = 10'b0;
assign pca_data_in_10b[1][19] = 10'b0;
assign pca_data_in_10b[1][20] = 10'b0;
assign pca_data_in_10b[1][21] = 10'b0;
assign pca_data_in_10b[1][22] = 10'b0;
assign pca_data_in_10b[1][23] = 10'b0;
assign pca_data_in_10b[1][24] = 10'b0;
assign pca_data_in_10b[1][25] = 10'b0;
assign pca_data_in_10b[1][26] = 10'b0;
assign pca_data_in_10b[1][27] = 10'b0;
assign pca_data_in_10b[1][28] = 10'b0;
assign pca_data_in_10b[1][29] = 10'b0;
assign pca_data_in_10b[1][30] = 10'b0;
assign pca_data_in_10b[1][31] = 10'b0;

// row 2 pixels 0-31 
assign pca_data_in_10b[2][0] = 10'b0;
assign pca_data_in_10b[2][1] = 10'b0;
assign pca_data_in_10b[2][2] = 10'b0;
assign pca_data_in_10b[2][3] = 10'b0;
assign pca_data_in_10b[2][4] = 10'b0;
assign pca_data_in_10b[2][5] = 10'b0;
assign pca_data_in_10b[2][6] = 10'b0;
assign pca_data_in_10b[2][7] = 10'b0;
assign pca_data_in_10b[2][8] = 10'b0;
assign pca_data_in_10b[2][9] = 10'b0;
assign pca_data_in_10b[2][10] = 10'b0;
assign pca_data_in_10b[2][11] = 10'b0;
assign pca_data_in_10b[2][12] = 10'b0;
assign pca_data_in_10b[2][13] = 10'b0;
assign pca_data_in_10b[2][14] = 10'b0;
assign pca_data_in_10b[2][15] = 10'b0;
assign pca_data_in_10b[2][16] = 10'b0;
assign pca_data_in_10b[2][17] = 10'b0;
assign pca_data_in_10b[2][18] = 10'b0;
assign pca_data_in_10b[2][19] = 10'b0;
assign pca_data_in_10b[2][20] = 10'b0;
assign pca_data_in_10b[2][21] = 10'b0;
assign pca_data_in_10b[2][22] = 10'b0;
assign pca_data_in_10b[2][23] = 10'b0;
assign pca_data_in_10b[2][24] = 10'b0;
assign pca_data_in_10b[2][25] = 10'b0;
assign pca_data_in_10b[2][26] = 10'b0;
assign pca_data_in_10b[2][27] = 10'b0;
assign pca_data_in_10b[2][28] = 10'b0;
assign pca_data_in_10b[2][29] = 10'b0;
assign pca_data_in_10b[2][30] = 10'b0;
assign pca_data_in_10b[2][31] = 10'b0;

// row 3 pixels 0-31 
assign pca_data_in_10b[3][0] = 10'b0;
assign pca_data_in_10b[3][1] = 10'b0;
assign pca_data_in_10b[3][2] = 10'b0;
assign pca_data_in_10b[3][3] = 10'b0;
assign pca_data_in_10b[3][4] = 10'b0;
assign pca_data_in_10b[3][5] = 10'b0;
assign pca_data_in_10b[3][6] = 10'b0;
assign pca_data_in_10b[3][7] = 10'b0;
assign pca_data_in_10b[3][8] = 10'b0;
assign pca_data_in_10b[3][9] = 10'b0;
assign pca_data_in_10b[3][10] = 10'b0;
assign pca_data_in_10b[3][11] = 10'b0;
assign pca_data_in_10b[3][12] = 10'b0;
assign pca_data_in_10b[3][13] = 10'b0;
assign pca_data_in_10b[3][14] = 10'b0;
assign pca_data_in_10b[3][15] = 10'b0;
assign pca_data_in_10b[3][16] = 10'b0;
assign pca_data_in_10b[3][17] = 10'b0;
assign pca_data_in_10b[3][18] = 10'b0;
assign pca_data_in_10b[3][19] = 10'b0;
assign pca_data_in_10b[3][20] = 10'b0;
assign pca_data_in_10b[3][21] = 10'b0;
assign pca_data_in_10b[3][22] = 10'b0;
assign pca_data_in_10b[3][23] = 10'b0;
assign pca_data_in_10b[3][24] = 10'b0;
assign pca_data_in_10b[3][25] = 10'b0;
assign pca_data_in_10b[3][26] = 10'b0;
assign pca_data_in_10b[3][27] = 10'b0;
assign pca_data_in_10b[3][28] = 10'b0;
assign pca_data_in_10b[3][29] = 10'b0;
assign pca_data_in_10b[3][30] = 10'b0;
assign pca_data_in_10b[3][31] = 10'b0;

// row 4 pixels 0-31 
assign pca_data_in_10b[4][0] = 10'b0;
assign pca_data_in_10b[4][1] = 10'b0;
assign pca_data_in_10b[4][2] = 10'b0;
assign pca_data_in_10b[4][3] = 10'b0;
assign pca_data_in_10b[4][4] = 10'b0;
assign pca_data_in_10b[4][5] = 10'b0;
assign pca_data_in_10b[4][6] = 10'b0;
assign pca_data_in_10b[4][7] = 10'b0;
assign pca_data_in_10b[4][8] = 10'b0;
assign pca_data_in_10b[4][9] = 10'b0;
assign pca_data_in_10b[4][10] = 10'b0;
assign pca_data_in_10b[4][11] = 10'b0;
assign pca_data_in_10b[4][12] = 10'b0;
assign pca_data_in_10b[4][13] = 10'b0;
assign pca_data_in_10b[4][14] = 10'b0;
assign pca_data_in_10b[4][15] = 10'b0;
assign pca_data_in_10b[4][16] = 10'b0;
assign pca_data_in_10b[4][17] = 10'b0;
assign pca_data_in_10b[4][18] = 10'b0;
assign pca_data_in_10b[4][19] = 10'b0;
assign pca_data_in_10b[4][20] = 10'b0;
assign pca_data_in_10b[4][21] = 10'b0;
assign pca_data_in_10b[4][22] = 10'b0;
assign pca_data_in_10b[4][23] = 10'b0;
assign pca_data_in_10b[4][24] = 10'b0;
assign pca_data_in_10b[4][25] = 10'b0;
assign pca_data_in_10b[4][26] = 10'b0;
assign pca_data_in_10b[4][27] = 10'b0;
assign pca_data_in_10b[4][28] = 10'b0;
assign pca_data_in_10b[4][29] = 10'b0;
assign pca_data_in_10b[4][30] = 10'b0;
assign pca_data_in_10b[4][31] = 10'b0;

// row 5 pixels 0-31 
assign pca_data_in_10b[5][0] = 10'b0;
assign pca_data_in_10b[5][1] = 10'b0;
assign pca_data_in_10b[5][2] = 10'b0;
assign pca_data_in_10b[5][3] = 10'b0;
assign pca_data_in_10b[5][4] = 10'b0;
assign pca_data_in_10b[5][5] = 10'b0;
assign pca_data_in_10b[5][6] = 10'b0;
assign pca_data_in_10b[5][7] = 10'b0;
assign pca_data_in_10b[5][8] = 10'b0;
assign pca_data_in_10b[5][9] = 10'b0;
assign pca_data_in_10b[5][10] = 10'b0;
assign pca_data_in_10b[5][11] = 10'b0;
assign pca_data_in_10b[5][12] = 10'b0;
assign pca_data_in_10b[5][13] = 10'b0;
assign pca_data_in_10b[5][14] = 10'b0;
assign pca_data_in_10b[5][15] = 10'b0;
assign pca_data_in_10b[5][16] = 10'b0;
assign pca_data_in_10b[5][17] = 10'b0;
assign pca_data_in_10b[5][18] = 10'b0;
assign pca_data_in_10b[5][19] = 10'b0;
assign pca_data_in_10b[5][20] = 10'b0;
assign pca_data_in_10b[5][21] = 10'b0;
assign pca_data_in_10b[5][22] = 10'b0;
assign pca_data_in_10b[5][23] = 10'b0;
assign pca_data_in_10b[5][24] = 10'b0;
assign pca_data_in_10b[5][25] = 10'b0;
assign pca_data_in_10b[5][26] = 10'b0;
assign pca_data_in_10b[5][27] = 10'b0;
assign pca_data_in_10b[5][28] = 10'b0;
assign pca_data_in_10b[5][29] = 10'b0;
assign pca_data_in_10b[5][30] = 10'b0;
assign pca_data_in_10b[5][31] = 10'b0;

// row 6 pixels 0-31 
assign pca_data_in_10b[6][0] = 10'b0;
assign pca_data_in_10b[6][1] = 10'b0;
assign pca_data_in_10b[6][2] = 10'b0;
assign pca_data_in_10b[6][3] = 10'b0;
assign pca_data_in_10b[6][4] = 10'b0;
assign pca_data_in_10b[6][5] = 10'b0;
assign pca_data_in_10b[6][6] = 10'b0;
assign pca_data_in_10b[6][7] = 10'b0;
assign pca_data_in_10b[6][8] = 10'b0;
assign pca_data_in_10b[6][9] = 10'b0;
assign pca_data_in_10b[6][10] = 10'b0;
assign pca_data_in_10b[6][11] = 10'b0;
assign pca_data_in_10b[6][12] = 10'b0;
assign pca_data_in_10b[6][13] = 10'b0;
assign pca_data_in_10b[6][14] = 10'b0;
assign pca_data_in_10b[6][15] = 10'b0;
assign pca_data_in_10b[6][16] = 10'b0;
assign pca_data_in_10b[6][17] = 10'b0;
assign pca_data_in_10b[6][18] = 10'b0;
assign pca_data_in_10b[6][19] = 10'b0;
assign pca_data_in_10b[6][20] = 10'b0;
assign pca_data_in_10b[6][21] = 10'b0;
assign pca_data_in_10b[6][22] = 10'b0;
assign pca_data_in_10b[6][23] = 10'b0;
assign pca_data_in_10b[6][24] = 10'b0;
assign pca_data_in_10b[6][25] = 10'b0;
assign pca_data_in_10b[6][26] = 10'b0;
assign pca_data_in_10b[6][27] = 10'b0;
assign pca_data_in_10b[6][28] = 10'b0;
assign pca_data_in_10b[6][29] = 10'b0;
assign pca_data_in_10b[6][30] = 10'b0;
assign pca_data_in_10b[6][31] = 10'b0;

// row 7 pixels 0-31 
assign pca_data_in_10b[7][0] = 10'b0;
assign pca_data_in_10b[7][1] = 10'b0;
assign pca_data_in_10b[7][2] = 10'b0;
assign pca_data_in_10b[7][3] = 10'b0;
assign pca_data_in_10b[7][4] = 10'b0;
assign pca_data_in_10b[7][5] = 10'b0;
assign pca_data_in_10b[7][6] = 10'b0;
assign pca_data_in_10b[7][7] = 10'b0;
assign pca_data_in_10b[7][8] = 10'b0;
assign pca_data_in_10b[7][9] = 10'b0;
assign pca_data_in_10b[7][10] = 10'b0;
assign pca_data_in_10b[7][11] = 10'b0;
assign pca_data_in_10b[7][12] = 10'b0;
assign pca_data_in_10b[7][13] = 10'b0;
assign pca_data_in_10b[7][14] = 10'b0;
assign pca_data_in_10b[7][15] = 10'b0;
assign pca_data_in_10b[7][16] = 10'b0;
assign pca_data_in_10b[7][17] = 10'b0;
assign pca_data_in_10b[7][18] = 10'b0;
assign pca_data_in_10b[7][19] = 10'b0;
assign pca_data_in_10b[7][20] = 10'b0;
assign pca_data_in_10b[7][21] = 10'b0;
assign pca_data_in_10b[7][22] = 10'b0;
assign pca_data_in_10b[7][23] = 10'b0;
assign pca_data_in_10b[7][24] = 10'b0;
assign pca_data_in_10b[7][25] = 10'b0;
assign pca_data_in_10b[7][26] = 10'b0;
assign pca_data_in_10b[7][27] = 10'b0;
assign pca_data_in_10b[7][28] = 10'b0;
assign pca_data_in_10b[7][29] = 10'b0;
assign pca_data_in_10b[7][30] = 10'b0;
assign pca_data_in_10b[7][31] = 10'b0;

// row 8 pixels 0-31 
assign pca_data_in_10b[8][0] = 10'b0;
assign pca_data_in_10b[8][1] = 10'b0;
assign pca_data_in_10b[8][2] = 10'b0;
assign pca_data_in_10b[8][3] = 10'b0;
assign pca_data_in_10b[8][4] = 10'b0;
assign pca_data_in_10b[8][5] = 10'b0;
assign pca_data_in_10b[8][6] = 10'b0;
assign pca_data_in_10b[8][7] = 10'b0;
assign pca_data_in_10b[8][8] = 10'b0;
assign pca_data_in_10b[8][9] = 10'b0;
assign pca_data_in_10b[8][10] = 10'b0;
assign pca_data_in_10b[8][11] = 10'b0;
assign pca_data_in_10b[8][12] = 10'b0;
assign pca_data_in_10b[8][13] = 10'b0;
assign pca_data_in_10b[8][14] = 10'b0;
assign pca_data_in_10b[8][15] = 10'b0;
assign pca_data_in_10b[8][16] = 10'b0;
assign pca_data_in_10b[8][17] = 10'b0;
assign pca_data_in_10b[8][18] = 10'b0;
assign pca_data_in_10b[8][19] = 10'b0;
assign pca_data_in_10b[8][20] = 10'b0;
assign pca_data_in_10b[8][21] = 10'b0;
assign pca_data_in_10b[8][22] = 10'b0;
assign pca_data_in_10b[8][23] = 10'b0;
assign pca_data_in_10b[8][24] = 10'b0;
assign pca_data_in_10b[8][25] = 10'b0;
assign pca_data_in_10b[8][26] = 10'b0;
assign pca_data_in_10b[8][27] = 10'b0;
assign pca_data_in_10b[8][28] = 10'b0;
assign pca_data_in_10b[8][29] = 10'b0;
assign pca_data_in_10b[8][30] = 10'b0;
assign pca_data_in_10b[8][31] = 10'b0;

// row 9 pixels 0-31 
assign pca_data_in_10b[9][0] = 10'b0;
assign pca_data_in_10b[9][1] = 10'b0;
assign pca_data_in_10b[9][2] = 10'b0;
assign pca_data_in_10b[9][3] = 10'b0;
assign pca_data_in_10b[9][4] = 10'b0;
assign pca_data_in_10b[9][5] = 10'b0;
assign pca_data_in_10b[9][6] = 10'b0;
assign pca_data_in_10b[9][7] = 10'b0;
assign pca_data_in_10b[9][8] = 10'b0;
assign pca_data_in_10b[9][9] = 10'b0;
assign pca_data_in_10b[9][10] = 10'b0;
assign pca_data_in_10b[9][11] = 10'b0;
assign pca_data_in_10b[9][12] = 10'b0;
assign pca_data_in_10b[9][13] = 10'b0;
assign pca_data_in_10b[9][14] = 10'b0;
assign pca_data_in_10b[9][15] = 10'b0;
assign pca_data_in_10b[9][16] = 10'b0;
assign pca_data_in_10b[9][17] = 10'b0;
assign pca_data_in_10b[9][18] = 10'b0;
assign pca_data_in_10b[9][19] = 10'b0;
assign pca_data_in_10b[9][20] = 10'b0;
assign pca_data_in_10b[9][21] = 10'b0;
assign pca_data_in_10b[9][22] = 10'b0;
assign pca_data_in_10b[9][23] = 10'b0;
assign pca_data_in_10b[9][24] = 10'b0;
assign pca_data_in_10b[9][25] = 10'b0;
assign pca_data_in_10b[9][26] = 10'b0;
assign pca_data_in_10b[9][27] = 10'b0;
assign pca_data_in_10b[9][28] = 10'b0;
assign pca_data_in_10b[9][29] = 10'b0;
assign pca_data_in_10b[9][30] = 10'b0;
assign pca_data_in_10b[9][31] = 10'b0;

// row 10 pixels 0-31 
assign pca_data_in_10b[10][0] = 10'b0;
assign pca_data_in_10b[10][1] = 10'b0;
assign pca_data_in_10b[10][2] = 10'b0;
assign pca_data_in_10b[10][3] = 10'b0;
assign pca_data_in_10b[10][4] = 10'b0;
assign pca_data_in_10b[10][5] = 10'b0;
assign pca_data_in_10b[10][6] = 10'b0;
assign pca_data_in_10b[10][7] = 10'b0;
assign pca_data_in_10b[10][8] = 10'b0;
assign pca_data_in_10b[10][9] = 10'b0;
assign pca_data_in_10b[10][10] = 10'b0;
assign pca_data_in_10b[10][11] = 10'b0;
assign pca_data_in_10b[10][12] = 10'b0;
assign pca_data_in_10b[10][13] = 10'b0;
assign pca_data_in_10b[10][14] = 10'b0;
assign pca_data_in_10b[10][15] = 10'b0;
assign pca_data_in_10b[10][16] = 10'b0;
assign pca_data_in_10b[10][17] = 10'b0;
assign pca_data_in_10b[10][18] = 10'b0;
assign pca_data_in_10b[10][19] = 10'b0;
assign pca_data_in_10b[10][20] = 10'b0;
assign pca_data_in_10b[10][21] = 10'b0;
assign pca_data_in_10b[10][22] = 10'b0;
assign pca_data_in_10b[10][23] = 10'b0;
assign pca_data_in_10b[10][24] = 10'b0;
assign pca_data_in_10b[10][25] = 10'b0;
assign pca_data_in_10b[10][26] = 10'b0;
assign pca_data_in_10b[10][27] = 10'b0;
assign pca_data_in_10b[10][28] = 10'b0;
assign pca_data_in_10b[10][29] = 10'b0;
assign pca_data_in_10b[10][30] = 10'b0;
assign pca_data_in_10b[10][31] = 10'b0;

// row 11 pixels 0-31 
assign pca_data_in_10b[11][0] = 10'b0;
assign pca_data_in_10b[11][1] = 10'b0;
assign pca_data_in_10b[11][2] = 10'b0;
assign pca_data_in_10b[11][3] = 10'b0;
assign pca_data_in_10b[11][4] = 10'b0;
assign pca_data_in_10b[11][5] = 10'b0;
assign pca_data_in_10b[11][6] = 10'b0;
assign pca_data_in_10b[11][7] = 10'b0;
assign pca_data_in_10b[11][8] = 10'b0;
assign pca_data_in_10b[11][9] = 10'b0;
assign pca_data_in_10b[11][10] = 10'b0;
assign pca_data_in_10b[11][11] = 10'b0;
assign pca_data_in_10b[11][12] = 10'b0;
assign pca_data_in_10b[11][13] = 10'b0;
assign pca_data_in_10b[11][14] = 10'b0;
assign pca_data_in_10b[11][15] = 10'b0;
assign pca_data_in_10b[11][16] = 10'b0;
assign pca_data_in_10b[11][17] = 10'b0;
assign pca_data_in_10b[11][18] = 10'b0;
assign pca_data_in_10b[11][19] = 10'b0;
assign pca_data_in_10b[11][20] = 10'b0;
assign pca_data_in_10b[11][21] = 10'b0;
assign pca_data_in_10b[11][22] = 10'b0;
assign pca_data_in_10b[11][23] = 10'b0;
assign pca_data_in_10b[11][24] = 10'b0;
assign pca_data_in_10b[11][25] = 10'b0;
assign pca_data_in_10b[11][26] = 10'b0;
assign pca_data_in_10b[11][27] = 10'b0;
assign pca_data_in_10b[11][28] = 10'b0;
assign pca_data_in_10b[11][29] = 10'b0;
assign pca_data_in_10b[11][30] = 10'b0;
assign pca_data_in_10b[11][31] = 10'b0;

// row 12 pixels 0-31 
assign pca_data_in_10b[12][0] = 10'b0;
assign pca_data_in_10b[12][1] = 10'b0;
assign pca_data_in_10b[12][2] = 10'b0;
assign pca_data_in_10b[12][3] = 10'b0;
assign pca_data_in_10b[12][4] = 10'b0;
assign pca_data_in_10b[12][5] = 10'b0;
assign pca_data_in_10b[12][6] = 10'b0;
assign pca_data_in_10b[12][7] = 10'b0;
assign pca_data_in_10b[12][8] = 10'b0;
assign pca_data_in_10b[12][9] = 10'b0;
assign pca_data_in_10b[12][10] = 10'b0;
assign pca_data_in_10b[12][11] = 10'b0;
assign pca_data_in_10b[12][12] = 10'b0;
assign pca_data_in_10b[12][13] = 10'b0;
assign pca_data_in_10b[12][14] = 10'b0;
assign pca_data_in_10b[12][15] = 10'b0;
assign pca_data_in_10b[12][16] = 10'b1;
assign pca_data_in_10b[12][17] = 10'b1;
assign pca_data_in_10b[12][18] = 10'b0;
assign pca_data_in_10b[12][19] = 10'b0;
assign pca_data_in_10b[12][20] = 10'b0;
assign pca_data_in_10b[12][21] = 10'b0;
assign pca_data_in_10b[12][22] = 10'b0;
assign pca_data_in_10b[12][23] = 10'b0;
assign pca_data_in_10b[12][24] = 10'b0;
assign pca_data_in_10b[12][25] = 10'b0;
assign pca_data_in_10b[12][26] = 10'b0;
assign pca_data_in_10b[12][27] = 10'b0;
assign pca_data_in_10b[12][28] = 10'b0;
assign pca_data_in_10b[12][29] = 10'b0;
assign pca_data_in_10b[12][30] = 10'b0;
assign pca_data_in_10b[12][31] = 10'b0;

// row 13 pixels 0-31 
assign pca_data_in_10b[13][0] = 10'b0;
assign pca_data_in_10b[13][1] = 10'b0;
assign pca_data_in_10b[13][2] = 10'b0;
assign pca_data_in_10b[13][3] = 10'b0;
assign pca_data_in_10b[13][4] = 10'b0;
assign pca_data_in_10b[13][5] = 10'b0;
assign pca_data_in_10b[13][6] = 10'b0;
assign pca_data_in_10b[13][7] = 10'b0;
assign pca_data_in_10b[13][8] = 10'b0;
assign pca_data_in_10b[13][9] = 10'b0;
assign pca_data_in_10b[13][10] = 10'b0;
assign pca_data_in_10b[13][11] = 10'b0;
assign pca_data_in_10b[13][12] = 10'b0;
assign pca_data_in_10b[13][13] = 10'b1;
assign pca_data_in_10b[13][14] = 10'b0;
assign pca_data_in_10b[13][15] = 10'b111;
assign pca_data_in_10b[13][16] = 10'b1011;
assign pca_data_in_10b[13][17] = 10'b110;
assign pca_data_in_10b[13][18] = 10'b1;
assign pca_data_in_10b[13][19] = 10'b0;
assign pca_data_in_10b[13][20] = 10'b0;
assign pca_data_in_10b[13][21] = 10'b0;
assign pca_data_in_10b[13][22] = 10'b0;
assign pca_data_in_10b[13][23] = 10'b0;
assign pca_data_in_10b[13][24] = 10'b0;
assign pca_data_in_10b[13][25] = 10'b0;
assign pca_data_in_10b[13][26] = 10'b0;
assign pca_data_in_10b[13][27] = 10'b0;
assign pca_data_in_10b[13][28] = 10'b0;
assign pca_data_in_10b[13][29] = 10'b0;
assign pca_data_in_10b[13][30] = 10'b0;
assign pca_data_in_10b[13][31] = 10'b0;

// row 14 pixels 0-31 
assign pca_data_in_10b[14][0] = 10'b0;
assign pca_data_in_10b[14][1] = 10'b0;
assign pca_data_in_10b[14][2] = 10'b0;
assign pca_data_in_10b[14][3] = 10'b0;
assign pca_data_in_10b[14][4] = 10'b0;
assign pca_data_in_10b[14][5] = 10'b0;
assign pca_data_in_10b[14][6] = 10'b0;
assign pca_data_in_10b[14][7] = 10'b0;
assign pca_data_in_10b[14][8] = 10'b0;
assign pca_data_in_10b[14][9] = 10'b0;
assign pca_data_in_10b[14][10] = 10'b0;
assign pca_data_in_10b[14][11] = 10'b0;
assign pca_data_in_10b[14][12] = 10'b0;
assign pca_data_in_10b[14][13] = 10'b1;
assign pca_data_in_10b[14][14] = 10'b1001;
assign pca_data_in_10b[14][15] = 10'b11011;
assign pca_data_in_10b[14][16] = 10'b1100001;
assign pca_data_in_10b[14][17] = 10'b101001;
assign pca_data_in_10b[14][18] = 10'b1001;
assign pca_data_in_10b[14][19] = 10'b0;
assign pca_data_in_10b[14][20] = 10'b0;
assign pca_data_in_10b[14][21] = 10'b0;
assign pca_data_in_10b[14][22] = 10'b0;
assign pca_data_in_10b[14][23] = 10'b0;
assign pca_data_in_10b[14][24] = 10'b0;
assign pca_data_in_10b[14][25] = 10'b0;
assign pca_data_in_10b[14][26] = 10'b0;
assign pca_data_in_10b[14][27] = 10'b0;
assign pca_data_in_10b[14][28] = 10'b0;
assign pca_data_in_10b[14][29] = 10'b0;
assign pca_data_in_10b[14][30] = 10'b0;
assign pca_data_in_10b[14][31] = 10'b0;

// row 15 pixels 0-31 
assign pca_data_in_10b[15][0] = 10'b0;
assign pca_data_in_10b[15][1] = 10'b0;
assign pca_data_in_10b[15][2] = 10'b0;
assign pca_data_in_10b[15][3] = 10'b0;
assign pca_data_in_10b[15][4] = 10'b0;
assign pca_data_in_10b[15][5] = 10'b0;
assign pca_data_in_10b[15][6] = 10'b0;
assign pca_data_in_10b[15][7] = 10'b0;
assign pca_data_in_10b[15][8] = 10'b0;
assign pca_data_in_10b[15][9] = 10'b0;
assign pca_data_in_10b[15][10] = 10'b0;
assign pca_data_in_10b[15][11] = 10'b0;
assign pca_data_in_10b[15][12] = 10'b0;
assign pca_data_in_10b[15][13] = 10'b1;
assign pca_data_in_10b[15][14] = 10'b101110;
assign pca_data_in_10b[15][15] = 10'b11110010;
assign pca_data_in_10b[15][16] = 10'b111010010;
assign pca_data_in_10b[15][17] = 10'b100001111;
assign pca_data_in_10b[15][18] = 10'b101100;
assign pca_data_in_10b[15][19] = 10'b101;
assign pca_data_in_10b[15][20] = 10'b0;
assign pca_data_in_10b[15][21] = 10'b0;
assign pca_data_in_10b[15][22] = 10'b0;
assign pca_data_in_10b[15][23] = 10'b0;
assign pca_data_in_10b[15][24] = 10'b0;
assign pca_data_in_10b[15][25] = 10'b0;
assign pca_data_in_10b[15][26] = 10'b0;
assign pca_data_in_10b[15][27] = 10'b0;
assign pca_data_in_10b[15][28] = 10'b0;
assign pca_data_in_10b[15][29] = 10'b0;
assign pca_data_in_10b[15][30] = 10'b0;
assign pca_data_in_10b[15][31] = 10'b0;

// row 16 pixels 0-31 
assign pca_data_in_10b[16][0] = 10'b0;
assign pca_data_in_10b[16][1] = 10'b0;
assign pca_data_in_10b[16][2] = 10'b0;
assign pca_data_in_10b[16][3] = 10'b0;
assign pca_data_in_10b[16][4] = 10'b0;
assign pca_data_in_10b[16][5] = 10'b0;
assign pca_data_in_10b[16][6] = 10'b0;
assign pca_data_in_10b[16][7] = 10'b0;
assign pca_data_in_10b[16][8] = 10'b0;
assign pca_data_in_10b[16][9] = 10'b0;
assign pca_data_in_10b[16][10] = 10'b0;
assign pca_data_in_10b[16][11] = 10'b0;
assign pca_data_in_10b[16][12] = 10'b1;
assign pca_data_in_10b[16][13] = 10'b100;
assign pca_data_in_10b[16][14] = 10'b1011000;
assign pca_data_in_10b[16][15] = 10'b111010010;
assign pca_data_in_10b[16][16] = 10'b1101001000;
assign pca_data_in_10b[16][17] = 10'b111010000;
assign pca_data_in_10b[16][18] = 10'b1011001;
assign pca_data_in_10b[16][19] = 10'b111;
assign pca_data_in_10b[16][20] = 10'b0;
assign pca_data_in_10b[16][21] = 10'b0;
assign pca_data_in_10b[16][22] = 10'b0;
assign pca_data_in_10b[16][23] = 10'b0;
assign pca_data_in_10b[16][24] = 10'b0;
assign pca_data_in_10b[16][25] = 10'b0;
assign pca_data_in_10b[16][26] = 10'b0;
assign pca_data_in_10b[16][27] = 10'b0;
assign pca_data_in_10b[16][28] = 10'b0;
assign pca_data_in_10b[16][29] = 10'b0;
assign pca_data_in_10b[16][30] = 10'b0;
assign pca_data_in_10b[16][31] = 10'b0;

// row 17 pixels 0-31 
assign pca_data_in_10b[17][0] = 10'b0;
assign pca_data_in_10b[17][1] = 10'b0;
assign pca_data_in_10b[17][2] = 10'b0;
assign pca_data_in_10b[17][3] = 10'b0;
assign pca_data_in_10b[17][4] = 10'b0;
assign pca_data_in_10b[17][5] = 10'b0;
assign pca_data_in_10b[17][6] = 10'b0;
assign pca_data_in_10b[17][7] = 10'b0;
assign pca_data_in_10b[17][8] = 10'b0;
assign pca_data_in_10b[17][9] = 10'b0;
assign pca_data_in_10b[17][10] = 10'b0;
assign pca_data_in_10b[17][11] = 10'b0;
assign pca_data_in_10b[17][12] = 10'b0;
assign pca_data_in_10b[17][13] = 10'b10;
assign pca_data_in_10b[17][14] = 10'b100101;
assign pca_data_in_10b[17][15] = 10'b11110100;
assign pca_data_in_10b[17][16] = 10'b111001011;
assign pca_data_in_10b[17][17] = 10'b100000000;
assign pca_data_in_10b[17][18] = 10'b101001;
assign pca_data_in_10b[17][19] = 10'b10;
assign pca_data_in_10b[17][20] = 10'b0;
assign pca_data_in_10b[17][21] = 10'b0;
assign pca_data_in_10b[17][22] = 10'b0;
assign pca_data_in_10b[17][23] = 10'b0;
assign pca_data_in_10b[17][24] = 10'b0;
assign pca_data_in_10b[17][25] = 10'b0;
assign pca_data_in_10b[17][26] = 10'b0;
assign pca_data_in_10b[17][27] = 10'b0;
assign pca_data_in_10b[17][28] = 10'b0;
assign pca_data_in_10b[17][29] = 10'b0;
assign pca_data_in_10b[17][30] = 10'b0;
assign pca_data_in_10b[17][31] = 10'b0;

// row 18 pixels 0-31 
assign pca_data_in_10b[18][0] = 10'b0;
assign pca_data_in_10b[18][1] = 10'b0;
assign pca_data_in_10b[18][2] = 10'b0;
assign pca_data_in_10b[18][3] = 10'b0;
assign pca_data_in_10b[18][4] = 10'b0;
assign pca_data_in_10b[18][5] = 10'b0;
assign pca_data_in_10b[18][6] = 10'b0;
assign pca_data_in_10b[18][7] = 10'b0;
assign pca_data_in_10b[18][8] = 10'b0;
assign pca_data_in_10b[18][9] = 10'b0;
assign pca_data_in_10b[18][10] = 10'b0;
assign pca_data_in_10b[18][11] = 10'b0;
assign pca_data_in_10b[18][12] = 10'b0;
assign pca_data_in_10b[18][13] = 10'b10;
assign pca_data_in_10b[18][14] = 10'b1011;
assign pca_data_in_10b[18][15] = 10'b101110;
assign pca_data_in_10b[18][16] = 10'b1010011;
assign pca_data_in_10b[18][17] = 10'b100111;
assign pca_data_in_10b[18][18] = 10'b1000;
assign pca_data_in_10b[18][19] = 10'b1;
assign pca_data_in_10b[18][20] = 10'b0;
assign pca_data_in_10b[18][21] = 10'b0;
assign pca_data_in_10b[18][22] = 10'b0;
assign pca_data_in_10b[18][23] = 10'b0;
assign pca_data_in_10b[18][24] = 10'b0;
assign pca_data_in_10b[18][25] = 10'b0;
assign pca_data_in_10b[18][26] = 10'b0;
assign pca_data_in_10b[18][27] = 10'b0;
assign pca_data_in_10b[18][28] = 10'b0;
assign pca_data_in_10b[18][29] = 10'b0;
assign pca_data_in_10b[18][30] = 10'b0;
assign pca_data_in_10b[18][31] = 10'b0;

// row 19 pixels 0-31 
assign pca_data_in_10b[19][0] = 10'b0;
assign pca_data_in_10b[19][1] = 10'b0;
assign pca_data_in_10b[19][2] = 10'b0;
assign pca_data_in_10b[19][3] = 10'b0;
assign pca_data_in_10b[19][4] = 10'b0;
assign pca_data_in_10b[19][5] = 10'b0;
assign pca_data_in_10b[19][6] = 10'b0;
assign pca_data_in_10b[19][7] = 10'b0;
assign pca_data_in_10b[19][8] = 10'b0;
assign pca_data_in_10b[19][9] = 10'b0;
assign pca_data_in_10b[19][10] = 10'b0;
assign pca_data_in_10b[19][11] = 10'b0;
assign pca_data_in_10b[19][12] = 10'b0;
assign pca_data_in_10b[19][13] = 10'b0;
assign pca_data_in_10b[19][14] = 10'b0;
assign pca_data_in_10b[19][15] = 10'b11;
assign pca_data_in_10b[19][16] = 10'b11;
assign pca_data_in_10b[19][17] = 10'b10;
assign pca_data_in_10b[19][18] = 10'b0;
assign pca_data_in_10b[19][19] = 10'b0;
assign pca_data_in_10b[19][20] = 10'b0;
assign pca_data_in_10b[19][21] = 10'b0;
assign pca_data_in_10b[19][22] = 10'b0;
assign pca_data_in_10b[19][23] = 10'b0;
assign pca_data_in_10b[19][24] = 10'b0;
assign pca_data_in_10b[19][25] = 10'b0;
assign pca_data_in_10b[19][26] = 10'b0;
assign pca_data_in_10b[19][27] = 10'b0;
assign pca_data_in_10b[19][28] = 10'b0;
assign pca_data_in_10b[19][29] = 10'b0;
assign pca_data_in_10b[19][30] = 10'b0;
assign pca_data_in_10b[19][31] = 10'b0;

// row 20 pixels 0-31 
assign pca_data_in_10b[20][0] = 10'b0;
assign pca_data_in_10b[20][1] = 10'b0;
assign pca_data_in_10b[20][2] = 10'b0;
assign pca_data_in_10b[20][3] = 10'b0;
assign pca_data_in_10b[20][4] = 10'b0;
assign pca_data_in_10b[20][5] = 10'b0;
assign pca_data_in_10b[20][6] = 10'b0;
assign pca_data_in_10b[20][7] = 10'b0;
assign pca_data_in_10b[20][8] = 10'b0;
assign pca_data_in_10b[20][9] = 10'b0;
assign pca_data_in_10b[20][10] = 10'b0;
assign pca_data_in_10b[20][11] = 10'b0;
assign pca_data_in_10b[20][12] = 10'b0;
assign pca_data_in_10b[20][13] = 10'b0;
assign pca_data_in_10b[20][14] = 10'b1;
assign pca_data_in_10b[20][15] = 10'b0;
assign pca_data_in_10b[20][16] = 10'b1;
assign pca_data_in_10b[20][17] = 10'b0;
assign pca_data_in_10b[20][18] = 10'b0;
assign pca_data_in_10b[20][19] = 10'b0;
assign pca_data_in_10b[20][20] = 10'b0;
assign pca_data_in_10b[20][21] = 10'b0;
assign pca_data_in_10b[20][22] = 10'b0;
assign pca_data_in_10b[20][23] = 10'b0;
assign pca_data_in_10b[20][24] = 10'b0;
assign pca_data_in_10b[20][25] = 10'b0;
assign pca_data_in_10b[20][26] = 10'b0;
assign pca_data_in_10b[20][27] = 10'b0;
assign pca_data_in_10b[20][28] = 10'b0;
assign pca_data_in_10b[20][29] = 10'b0;
assign pca_data_in_10b[20][30] = 10'b0;
assign pca_data_in_10b[20][31] = 10'b0;

// row 21 pixels 0-31 
assign pca_data_in_10b[21][0] = 10'b0;
assign pca_data_in_10b[21][1] = 10'b0;
assign pca_data_in_10b[21][2] = 10'b0;
assign pca_data_in_10b[21][3] = 10'b0;
assign pca_data_in_10b[21][4] = 10'b0;
assign pca_data_in_10b[21][5] = 10'b0;
assign pca_data_in_10b[21][6] = 10'b0;
assign pca_data_in_10b[21][7] = 10'b0;
assign pca_data_in_10b[21][8] = 10'b0;
assign pca_data_in_10b[21][9] = 10'b0;
assign pca_data_in_10b[21][10] = 10'b0;
assign pca_data_in_10b[21][11] = 10'b0;
assign pca_data_in_10b[21][12] = 10'b0;
assign pca_data_in_10b[21][13] = 10'b0;
assign pca_data_in_10b[21][14] = 10'b0;
assign pca_data_in_10b[21][15] = 10'b1;
assign pca_data_in_10b[21][16] = 10'b0;
assign pca_data_in_10b[21][17] = 10'b0;
assign pca_data_in_10b[21][18] = 10'b0;
assign pca_data_in_10b[21][19] = 10'b0;
assign pca_data_in_10b[21][20] = 10'b0;
assign pca_data_in_10b[21][21] = 10'b0;
assign pca_data_in_10b[21][22] = 10'b0;
assign pca_data_in_10b[21][23] = 10'b0;
assign pca_data_in_10b[21][24] = 10'b0;
assign pca_data_in_10b[21][25] = 10'b0;
assign pca_data_in_10b[21][26] = 10'b0;
assign pca_data_in_10b[21][27] = 10'b0;
assign pca_data_in_10b[21][28] = 10'b0;
assign pca_data_in_10b[21][29] = 10'b0;
assign pca_data_in_10b[21][30] = 10'b0;
assign pca_data_in_10b[21][31] = 10'b0;

// row 22 pixels 0-31 
assign pca_data_in_10b[22][0] = 10'b0;
assign pca_data_in_10b[22][1] = 10'b0;
assign pca_data_in_10b[22][2] = 10'b0;
assign pca_data_in_10b[22][3] = 10'b0;
assign pca_data_in_10b[22][4] = 10'b0;
assign pca_data_in_10b[22][5] = 10'b0;
assign pca_data_in_10b[22][6] = 10'b0;
assign pca_data_in_10b[22][7] = 10'b0;
assign pca_data_in_10b[22][8] = 10'b0;
assign pca_data_in_10b[22][9] = 10'b0;
assign pca_data_in_10b[22][10] = 10'b0;
assign pca_data_in_10b[22][11] = 10'b0;
assign pca_data_in_10b[22][12] = 10'b0;
assign pca_data_in_10b[22][13] = 10'b0;
assign pca_data_in_10b[22][14] = 10'b0;
assign pca_data_in_10b[22][15] = 10'b0;
assign pca_data_in_10b[22][16] = 10'b0;
assign pca_data_in_10b[22][17] = 10'b0;
assign pca_data_in_10b[22][18] = 10'b0;
assign pca_data_in_10b[22][19] = 10'b0;
assign pca_data_in_10b[22][20] = 10'b0;
assign pca_data_in_10b[22][21] = 10'b0;
assign pca_data_in_10b[22][22] = 10'b0;
assign pca_data_in_10b[22][23] = 10'b0;
assign pca_data_in_10b[22][24] = 10'b0;
assign pca_data_in_10b[22][25] = 10'b0;
assign pca_data_in_10b[22][26] = 10'b0;
assign pca_data_in_10b[22][27] = 10'b0;
assign pca_data_in_10b[22][28] = 10'b0;
assign pca_data_in_10b[22][29] = 10'b0;
assign pca_data_in_10b[22][30] = 10'b0;
assign pca_data_in_10b[22][31] = 10'b0;

// row 23 pixels 0-31 
assign pca_data_in_10b[23][0] = 10'b0;
assign pca_data_in_10b[23][1] = 10'b0;
assign pca_data_in_10b[23][2] = 10'b0;
assign pca_data_in_10b[23][3] = 10'b0;
assign pca_data_in_10b[23][4] = 10'b0;
assign pca_data_in_10b[23][5] = 10'b0;
assign pca_data_in_10b[23][6] = 10'b0;
assign pca_data_in_10b[23][7] = 10'b0;
assign pca_data_in_10b[23][8] = 10'b0;
assign pca_data_in_10b[23][9] = 10'b0;
assign pca_data_in_10b[23][10] = 10'b0;
assign pca_data_in_10b[23][11] = 10'b0;
assign pca_data_in_10b[23][12] = 10'b0;
assign pca_data_in_10b[23][13] = 10'b0;
assign pca_data_in_10b[23][14] = 10'b0;
assign pca_data_in_10b[23][15] = 10'b0;
assign pca_data_in_10b[23][16] = 10'b0;
assign pca_data_in_10b[23][17] = 10'b0;
assign pca_data_in_10b[23][18] = 10'b0;
assign pca_data_in_10b[23][19] = 10'b0;
assign pca_data_in_10b[23][20] = 10'b0;
assign pca_data_in_10b[23][21] = 10'b0;
assign pca_data_in_10b[23][22] = 10'b0;
assign pca_data_in_10b[23][23] = 10'b0;
assign pca_data_in_10b[23][24] = 10'b0;
assign pca_data_in_10b[23][25] = 10'b0;
assign pca_data_in_10b[23][26] = 10'b0;
assign pca_data_in_10b[23][27] = 10'b0;
assign pca_data_in_10b[23][28] = 10'b0;
assign pca_data_in_10b[23][29] = 10'b0;
assign pca_data_in_10b[23][30] = 10'b0;
assign pca_data_in_10b[23][31] = 10'b0;

// row 24 pixels 0-31 
assign pca_data_in_10b[24][0] = 10'b0;
assign pca_data_in_10b[24][1] = 10'b0;
assign pca_data_in_10b[24][2] = 10'b0;
assign pca_data_in_10b[24][3] = 10'b0;
assign pca_data_in_10b[24][4] = 10'b0;
assign pca_data_in_10b[24][5] = 10'b0;
assign pca_data_in_10b[24][6] = 10'b0;
assign pca_data_in_10b[24][7] = 10'b0;
assign pca_data_in_10b[24][8] = 10'b0;
assign pca_data_in_10b[24][9] = 10'b0;
assign pca_data_in_10b[24][10] = 10'b0;
assign pca_data_in_10b[24][11] = 10'b0;
assign pca_data_in_10b[24][12] = 10'b0;
assign pca_data_in_10b[24][13] = 10'b0;
assign pca_data_in_10b[24][14] = 10'b0;
assign pca_data_in_10b[24][15] = 10'b0;
assign pca_data_in_10b[24][16] = 10'b0;
assign pca_data_in_10b[24][17] = 10'b0;
assign pca_data_in_10b[24][18] = 10'b0;
assign pca_data_in_10b[24][19] = 10'b0;
assign pca_data_in_10b[24][20] = 10'b0;
assign pca_data_in_10b[24][21] = 10'b0;
assign pca_data_in_10b[24][22] = 10'b0;
assign pca_data_in_10b[24][23] = 10'b0;
assign pca_data_in_10b[24][24] = 10'b0;
assign pca_data_in_10b[24][25] = 10'b0;
assign pca_data_in_10b[24][26] = 10'b0;
assign pca_data_in_10b[24][27] = 10'b0;
assign pca_data_in_10b[24][28] = 10'b0;
assign pca_data_in_10b[24][29] = 10'b0;
assign pca_data_in_10b[24][30] = 10'b0;
assign pca_data_in_10b[24][31] = 10'b0;

// row 25 pixels 0-31 
assign pca_data_in_10b[25][0] = 10'b0;
assign pca_data_in_10b[25][1] = 10'b0;
assign pca_data_in_10b[25][2] = 10'b0;
assign pca_data_in_10b[25][3] = 10'b0;
assign pca_data_in_10b[25][4] = 10'b0;
assign pca_data_in_10b[25][5] = 10'b0;
assign pca_data_in_10b[25][6] = 10'b0;
assign pca_data_in_10b[25][7] = 10'b0;
assign pca_data_in_10b[25][8] = 10'b0;
assign pca_data_in_10b[25][9] = 10'b0;
assign pca_data_in_10b[25][10] = 10'b0;
assign pca_data_in_10b[25][11] = 10'b0;
assign pca_data_in_10b[25][12] = 10'b0;
assign pca_data_in_10b[25][13] = 10'b0;
assign pca_data_in_10b[25][14] = 10'b0;
assign pca_data_in_10b[25][15] = 10'b0;
assign pca_data_in_10b[25][16] = 10'b0;
assign pca_data_in_10b[25][17] = 10'b0;
assign pca_data_in_10b[25][18] = 10'b0;
assign pca_data_in_10b[25][19] = 10'b0;
assign pca_data_in_10b[25][20] = 10'b0;
assign pca_data_in_10b[25][21] = 10'b0;
assign pca_data_in_10b[25][22] = 10'b0;
assign pca_data_in_10b[25][23] = 10'b0;
assign pca_data_in_10b[25][24] = 10'b0;
assign pca_data_in_10b[25][25] = 10'b0;
assign pca_data_in_10b[25][26] = 10'b0;
assign pca_data_in_10b[25][27] = 10'b0;
assign pca_data_in_10b[25][28] = 10'b0;
assign pca_data_in_10b[25][29] = 10'b0;
assign pca_data_in_10b[25][30] = 10'b0;
assign pca_data_in_10b[25][31] = 10'b0;

// row 26 pixels 0-31 
assign pca_data_in_10b[26][0] = 10'b0;
assign pca_data_in_10b[26][1] = 10'b0;
assign pca_data_in_10b[26][2] = 10'b0;
assign pca_data_in_10b[26][3] = 10'b0;
assign pca_data_in_10b[26][4] = 10'b0;
assign pca_data_in_10b[26][5] = 10'b0;
assign pca_data_in_10b[26][6] = 10'b0;
assign pca_data_in_10b[26][7] = 10'b0;
assign pca_data_in_10b[26][8] = 10'b0;
assign pca_data_in_10b[26][9] = 10'b0;
assign pca_data_in_10b[26][10] = 10'b0;
assign pca_data_in_10b[26][11] = 10'b0;
assign pca_data_in_10b[26][12] = 10'b0;
assign pca_data_in_10b[26][13] = 10'b0;
assign pca_data_in_10b[26][14] = 10'b0;
assign pca_data_in_10b[26][15] = 10'b0;
assign pca_data_in_10b[26][16] = 10'b0;
assign pca_data_in_10b[26][17] = 10'b0;
assign pca_data_in_10b[26][18] = 10'b0;
assign pca_data_in_10b[26][19] = 10'b0;
assign pca_data_in_10b[26][20] = 10'b0;
assign pca_data_in_10b[26][21] = 10'b0;
assign pca_data_in_10b[26][22] = 10'b0;
assign pca_data_in_10b[26][23] = 10'b0;
assign pca_data_in_10b[26][24] = 10'b0;
assign pca_data_in_10b[26][25] = 10'b0;
assign pca_data_in_10b[26][26] = 10'b0;
assign pca_data_in_10b[26][27] = 10'b0;
assign pca_data_in_10b[26][28] = 10'b0;
assign pca_data_in_10b[26][29] = 10'b0;
assign pca_data_in_10b[26][30] = 10'b0;
assign pca_data_in_10b[26][31] = 10'b0;

// row 27 pixels 0-31 
assign pca_data_in_10b[27][0] = 10'b0;
assign pca_data_in_10b[27][1] = 10'b0;
assign pca_data_in_10b[27][2] = 10'b0;
assign pca_data_in_10b[27][3] = 10'b0;
assign pca_data_in_10b[27][4] = 10'b0;
assign pca_data_in_10b[27][5] = 10'b0;
assign pca_data_in_10b[27][6] = 10'b0;
assign pca_data_in_10b[27][7] = 10'b0;
assign pca_data_in_10b[27][8] = 10'b0;
assign pca_data_in_10b[27][9] = 10'b0;
assign pca_data_in_10b[27][10] = 10'b0;
assign pca_data_in_10b[27][11] = 10'b0;
assign pca_data_in_10b[27][12] = 10'b0;
assign pca_data_in_10b[27][13] = 10'b0;
assign pca_data_in_10b[27][14] = 10'b0;
assign pca_data_in_10b[27][15] = 10'b0;
assign pca_data_in_10b[27][16] = 10'b0;
assign pca_data_in_10b[27][17] = 10'b0;
assign pca_data_in_10b[27][18] = 10'b0;
assign pca_data_in_10b[27][19] = 10'b0;
assign pca_data_in_10b[27][20] = 10'b0;
assign pca_data_in_10b[27][21] = 10'b0;
assign pca_data_in_10b[27][22] = 10'b0;
assign pca_data_in_10b[27][23] = 10'b0;
assign pca_data_in_10b[27][24] = 10'b0;
assign pca_data_in_10b[27][25] = 10'b0;
assign pca_data_in_10b[27][26] = 10'b0;
assign pca_data_in_10b[27][27] = 10'b0;
assign pca_data_in_10b[27][28] = 10'b0;
assign pca_data_in_10b[27][29] = 10'b0;
assign pca_data_in_10b[27][30] = 10'b0;
assign pca_data_in_10b[27][31] = 10'b0;

// row 28 pixels 0-31 
assign pca_data_in_10b[28][0] = 10'b0;
assign pca_data_in_10b[28][1] = 10'b0;
assign pca_data_in_10b[28][2] = 10'b0;
assign pca_data_in_10b[28][3] = 10'b0;
assign pca_data_in_10b[28][4] = 10'b0;
assign pca_data_in_10b[28][5] = 10'b0;
assign pca_data_in_10b[28][6] = 10'b0;
assign pca_data_in_10b[28][7] = 10'b0;
assign pca_data_in_10b[28][8] = 10'b0;
assign pca_data_in_10b[28][9] = 10'b0;
assign pca_data_in_10b[28][10] = 10'b0;
assign pca_data_in_10b[28][11] = 10'b0;
assign pca_data_in_10b[28][12] = 10'b0;
assign pca_data_in_10b[28][13] = 10'b0;
assign pca_data_in_10b[28][14] = 10'b0;
assign pca_data_in_10b[28][15] = 10'b0;
assign pca_data_in_10b[28][16] = 10'b0;
assign pca_data_in_10b[28][17] = 10'b0;
assign pca_data_in_10b[28][18] = 10'b0;
assign pca_data_in_10b[28][19] = 10'b0;
assign pca_data_in_10b[28][20] = 10'b0;
assign pca_data_in_10b[28][21] = 10'b0;
assign pca_data_in_10b[28][22] = 10'b0;
assign pca_data_in_10b[28][23] = 10'b0;
assign pca_data_in_10b[28][24] = 10'b0;
assign pca_data_in_10b[28][25] = 10'b0;
assign pca_data_in_10b[28][26] = 10'b0;
assign pca_data_in_10b[28][27] = 10'b0;
assign pca_data_in_10b[28][28] = 10'b0;
assign pca_data_in_10b[28][29] = 10'b0;
assign pca_data_in_10b[28][30] = 10'b0;
assign pca_data_in_10b[28][31] = 10'b0;

// row 29 pixels 0-31 
assign pca_data_in_10b[29][0] = 10'b0;
assign pca_data_in_10b[29][1] = 10'b0;
assign pca_data_in_10b[29][2] = 10'b0;
assign pca_data_in_10b[29][3] = 10'b0;
assign pca_data_in_10b[29][4] = 10'b0;
assign pca_data_in_10b[29][5] = 10'b0;
assign pca_data_in_10b[29][6] = 10'b0;
assign pca_data_in_10b[29][7] = 10'b0;
assign pca_data_in_10b[29][8] = 10'b0;
assign pca_data_in_10b[29][9] = 10'b0;
assign pca_data_in_10b[29][10] = 10'b0;
assign pca_data_in_10b[29][11] = 10'b0;
assign pca_data_in_10b[29][12] = 10'b0;
assign pca_data_in_10b[29][13] = 10'b0;
assign pca_data_in_10b[29][14] = 10'b0;
assign pca_data_in_10b[29][15] = 10'b0;
assign pca_data_in_10b[29][16] = 10'b0;
assign pca_data_in_10b[29][17] = 10'b0;
assign pca_data_in_10b[29][18] = 10'b0;
assign pca_data_in_10b[29][19] = 10'b0;
assign pca_data_in_10b[29][20] = 10'b0;
assign pca_data_in_10b[29][21] = 10'b0;
assign pca_data_in_10b[29][22] = 10'b0;
assign pca_data_in_10b[29][23] = 10'b0;
assign pca_data_in_10b[29][24] = 10'b0;
assign pca_data_in_10b[29][25] = 10'b0;
assign pca_data_in_10b[29][26] = 10'b0;
assign pca_data_in_10b[29][27] = 10'b0;
assign pca_data_in_10b[29][28] = 10'b0;
assign pca_data_in_10b[29][29] = 10'b0;
assign pca_data_in_10b[29][30] = 10'b0;
assign pca_data_in_10b[29][31] = 10'b0;

// row 30 pixels 0-31 
assign pca_data_in_10b[30][0] = 10'b0;
assign pca_data_in_10b[30][1] = 10'b0;
assign pca_data_in_10b[30][2] = 10'b0;
assign pca_data_in_10b[30][3] = 10'b0;
assign pca_data_in_10b[30][4] = 10'b0;
assign pca_data_in_10b[30][5] = 10'b0;
assign pca_data_in_10b[30][6] = 10'b0;
assign pca_data_in_10b[30][7] = 10'b0;
assign pca_data_in_10b[30][8] = 10'b0;
assign pca_data_in_10b[30][9] = 10'b0;
assign pca_data_in_10b[30][10] = 10'b0;
assign pca_data_in_10b[30][11] = 10'b0;
assign pca_data_in_10b[30][12] = 10'b0;
assign pca_data_in_10b[30][13] = 10'b0;
assign pca_data_in_10b[30][14] = 10'b0;
assign pca_data_in_10b[30][15] = 10'b0;
assign pca_data_in_10b[30][16] = 10'b0;
assign pca_data_in_10b[30][17] = 10'b0;
assign pca_data_in_10b[30][18] = 10'b0;
assign pca_data_in_10b[30][19] = 10'b0;
assign pca_data_in_10b[30][20] = 10'b0;
assign pca_data_in_10b[30][21] = 10'b0;
assign pca_data_in_10b[30][22] = 10'b0;
assign pca_data_in_10b[30][23] = 10'b0;
assign pca_data_in_10b[30][24] = 10'b0;
assign pca_data_in_10b[30][25] = 10'b0;
assign pca_data_in_10b[30][26] = 10'b0;
assign pca_data_in_10b[30][27] = 10'b0;
assign pca_data_in_10b[30][28] = 10'b0;
assign pca_data_in_10b[30][29] = 10'b0;
assign pca_data_in_10b[30][30] = 10'b0;
assign pca_data_in_10b[30][31] = 10'b0;

// row 31 pixels 0-31 
assign pca_data_in_10b[31][0] = 10'b0;
assign pca_data_in_10b[31][1] = 10'b0;
assign pca_data_in_10b[31][2] = 10'b0;
assign pca_data_in_10b[31][3] = 10'b0;
assign pca_data_in_10b[31][4] = 10'b0;
assign pca_data_in_10b[31][5] = 10'b0;
assign pca_data_in_10b[31][6] = 10'b0;
assign pca_data_in_10b[31][7] = 10'b0;
assign pca_data_in_10b[31][8] = 10'b0;
assign pca_data_in_10b[31][9] = 10'b0;
assign pca_data_in_10b[31][10] = 10'b0;
assign pca_data_in_10b[31][11] = 10'b0;
assign pca_data_in_10b[31][12] = 10'b0;
assign pca_data_in_10b[31][13] = 10'b0;
assign pca_data_in_10b[31][14] = 10'b0;
assign pca_data_in_10b[31][15] = 10'b0;
assign pca_data_in_10b[31][16] = 10'b0;
assign pca_data_in_10b[31][17] = 10'b0;
assign pca_data_in_10b[31][18] = 10'b0;
assign pca_data_in_10b[31][19] = 10'b0;
assign pca_data_in_10b[31][20] = 10'b0;
assign pca_data_in_10b[31][21] = 10'b0;
assign pca_data_in_10b[31][22] = 10'b0;
assign pca_data_in_10b[31][23] = 10'b0;
assign pca_data_in_10b[31][24] = 10'b0;
assign pca_data_in_10b[31][25] = 10'b0;
assign pca_data_in_10b[31][26] = 10'b0;
assign pca_data_in_10b[31][27] = 10'b0;
assign pca_data_in_10b[31][28] = 10'b0;
assign pca_data_in_10b[31][29] = 10'b0;
assign pca_data_in_10b[31][30] = 10'b0;
assign pca_data_in_10b[31][31] = 10'b0;


// 5b inputs to AE algorithm (after 3-range pseudo-log)


// row 0 pixels 0-31 
assign ae_data_in_5b[0][0] = 5'b0;
assign ae_data_in_5b[0][1] = 5'b0;
assign ae_data_in_5b[0][2] = 5'b0;
assign ae_data_in_5b[0][3] = 5'b0;
assign ae_data_in_5b[0][4] = 5'b0;
assign ae_data_in_5b[0][5] = 5'b0;
assign ae_data_in_5b[0][6] = 5'b0;
assign ae_data_in_5b[0][7] = 5'b0;
assign ae_data_in_5b[0][8] = 5'b0;
assign ae_data_in_5b[0][9] = 5'b0;
assign ae_data_in_5b[0][10] = 5'b0;
assign ae_data_in_5b[0][11] = 5'b0;
assign ae_data_in_5b[0][12] = 5'b0;
assign ae_data_in_5b[0][13] = 5'b0;
assign ae_data_in_5b[0][14] = 5'b0;
assign ae_data_in_5b[0][15] = 5'b0;
assign ae_data_in_5b[0][16] = 5'b0;
assign ae_data_in_5b[0][17] = 5'b0;
assign ae_data_in_5b[0][18] = 5'b0;
assign ae_data_in_5b[0][19] = 5'b0;
assign ae_data_in_5b[0][20] = 5'b0;
assign ae_data_in_5b[0][21] = 5'b0;
assign ae_data_in_5b[0][22] = 5'b0;
assign ae_data_in_5b[0][23] = 5'b0;
assign ae_data_in_5b[0][24] = 5'b0;
assign ae_data_in_5b[0][25] = 5'b0;
assign ae_data_in_5b[0][26] = 5'b0;
assign ae_data_in_5b[0][27] = 5'b0;
assign ae_data_in_5b[0][28] = 5'b0;
assign ae_data_in_5b[0][29] = 5'b0;
assign ae_data_in_5b[0][30] = 5'b0;
assign ae_data_in_5b[0][31] = 5'b0;

// row 1 pixels 0-31 
assign ae_data_in_5b[1][0] = 5'b0;
assign ae_data_in_5b[1][1] = 5'b0;
assign ae_data_in_5b[1][2] = 5'b0;
assign ae_data_in_5b[1][3] = 5'b0;
assign ae_data_in_5b[1][4] = 5'b0;
assign ae_data_in_5b[1][5] = 5'b0;
assign ae_data_in_5b[1][6] = 5'b0;
assign ae_data_in_5b[1][7] = 5'b0;
assign ae_data_in_5b[1][8] = 5'b0;
assign ae_data_in_5b[1][9] = 5'b0;
assign ae_data_in_5b[1][10] = 5'b0;
assign ae_data_in_5b[1][11] = 5'b0;
assign ae_data_in_5b[1][12] = 5'b0;
assign ae_data_in_5b[1][13] = 5'b0;
assign ae_data_in_5b[1][14] = 5'b0;
assign ae_data_in_5b[1][15] = 5'b0;
assign ae_data_in_5b[1][16] = 5'b0;
assign ae_data_in_5b[1][17] = 5'b0;
assign ae_data_in_5b[1][18] = 5'b0;
assign ae_data_in_5b[1][19] = 5'b0;
assign ae_data_in_5b[1][20] = 5'b0;
assign ae_data_in_5b[1][21] = 5'b0;
assign ae_data_in_5b[1][22] = 5'b0;
assign ae_data_in_5b[1][23] = 5'b0;
assign ae_data_in_5b[1][24] = 5'b0;
assign ae_data_in_5b[1][25] = 5'b0;
assign ae_data_in_5b[1][26] = 5'b0;
assign ae_data_in_5b[1][27] = 5'b0;
assign ae_data_in_5b[1][28] = 5'b0;
assign ae_data_in_5b[1][29] = 5'b0;
assign ae_data_in_5b[1][30] = 5'b0;
assign ae_data_in_5b[1][31] = 5'b0;

// row 2 pixels 0-31 
assign ae_data_in_5b[2][0] = 5'b0;
assign ae_data_in_5b[2][1] = 5'b0;
assign ae_data_in_5b[2][2] = 5'b0;
assign ae_data_in_5b[2][3] = 5'b0;
assign ae_data_in_5b[2][4] = 5'b0;
assign ae_data_in_5b[2][5] = 5'b0;
assign ae_data_in_5b[2][6] = 5'b0;
assign ae_data_in_5b[2][7] = 5'b0;
assign ae_data_in_5b[2][8] = 5'b0;
assign ae_data_in_5b[2][9] = 5'b0;
assign ae_data_in_5b[2][10] = 5'b0;
assign ae_data_in_5b[2][11] = 5'b0;
assign ae_data_in_5b[2][12] = 5'b0;
assign ae_data_in_5b[2][13] = 5'b0;
assign ae_data_in_5b[2][14] = 5'b0;
assign ae_data_in_5b[2][15] = 5'b0;
assign ae_data_in_5b[2][16] = 5'b0;
assign ae_data_in_5b[2][17] = 5'b0;
assign ae_data_in_5b[2][18] = 5'b0;
assign ae_data_in_5b[2][19] = 5'b0;
assign ae_data_in_5b[2][20] = 5'b0;
assign ae_data_in_5b[2][21] = 5'b0;
assign ae_data_in_5b[2][22] = 5'b0;
assign ae_data_in_5b[2][23] = 5'b0;
assign ae_data_in_5b[2][24] = 5'b0;
assign ae_data_in_5b[2][25] = 5'b0;
assign ae_data_in_5b[2][26] = 5'b0;
assign ae_data_in_5b[2][27] = 5'b0;
assign ae_data_in_5b[2][28] = 5'b0;
assign ae_data_in_5b[2][29] = 5'b0;
assign ae_data_in_5b[2][30] = 5'b0;
assign ae_data_in_5b[2][31] = 5'b0;

// row 3 pixels 0-31 
assign ae_data_in_5b[3][0] = 5'b0;
assign ae_data_in_5b[3][1] = 5'b0;
assign ae_data_in_5b[3][2] = 5'b0;
assign ae_data_in_5b[3][3] = 5'b0;
assign ae_data_in_5b[3][4] = 5'b0;
assign ae_data_in_5b[3][5] = 5'b0;
assign ae_data_in_5b[3][6] = 5'b0;
assign ae_data_in_5b[3][7] = 5'b0;
assign ae_data_in_5b[3][8] = 5'b0;
assign ae_data_in_5b[3][9] = 5'b0;
assign ae_data_in_5b[3][10] = 5'b0;
assign ae_data_in_5b[3][11] = 5'b0;
assign ae_data_in_5b[3][12] = 5'b0;
assign ae_data_in_5b[3][13] = 5'b0;
assign ae_data_in_5b[3][14] = 5'b0;
assign ae_data_in_5b[3][15] = 5'b0;
assign ae_data_in_5b[3][16] = 5'b0;
assign ae_data_in_5b[3][17] = 5'b0;
assign ae_data_in_5b[3][18] = 5'b0;
assign ae_data_in_5b[3][19] = 5'b0;
assign ae_data_in_5b[3][20] = 5'b0;
assign ae_data_in_5b[3][21] = 5'b0;
assign ae_data_in_5b[3][22] = 5'b0;
assign ae_data_in_5b[3][23] = 5'b0;
assign ae_data_in_5b[3][24] = 5'b0;
assign ae_data_in_5b[3][25] = 5'b0;
assign ae_data_in_5b[3][26] = 5'b0;
assign ae_data_in_5b[3][27] = 5'b0;
assign ae_data_in_5b[3][28] = 5'b0;
assign ae_data_in_5b[3][29] = 5'b0;
assign ae_data_in_5b[3][30] = 5'b0;
assign ae_data_in_5b[3][31] = 5'b0;

// row 4 pixels 0-31 
assign ae_data_in_5b[4][0] = 5'b0;
assign ae_data_in_5b[4][1] = 5'b0;
assign ae_data_in_5b[4][2] = 5'b0;
assign ae_data_in_5b[4][3] = 5'b0;
assign ae_data_in_5b[4][4] = 5'b0;
assign ae_data_in_5b[4][5] = 5'b0;
assign ae_data_in_5b[4][6] = 5'b0;
assign ae_data_in_5b[4][7] = 5'b0;
assign ae_data_in_5b[4][8] = 5'b0;
assign ae_data_in_5b[4][9] = 5'b0;
assign ae_data_in_5b[4][10] = 5'b0;
assign ae_data_in_5b[4][11] = 5'b0;
assign ae_data_in_5b[4][12] = 5'b0;
assign ae_data_in_5b[4][13] = 5'b0;
assign ae_data_in_5b[4][14] = 5'b0;
assign ae_data_in_5b[4][15] = 5'b0;
assign ae_data_in_5b[4][16] = 5'b0;
assign ae_data_in_5b[4][17] = 5'b0;
assign ae_data_in_5b[4][18] = 5'b0;
assign ae_data_in_5b[4][19] = 5'b0;
assign ae_data_in_5b[4][20] = 5'b0;
assign ae_data_in_5b[4][21] = 5'b0;
assign ae_data_in_5b[4][22] = 5'b0;
assign ae_data_in_5b[4][23] = 5'b0;
assign ae_data_in_5b[4][24] = 5'b0;
assign ae_data_in_5b[4][25] = 5'b0;
assign ae_data_in_5b[4][26] = 5'b0;
assign ae_data_in_5b[4][27] = 5'b0;
assign ae_data_in_5b[4][28] = 5'b0;
assign ae_data_in_5b[4][29] = 5'b0;
assign ae_data_in_5b[4][30] = 5'b0;
assign ae_data_in_5b[4][31] = 5'b0;

// row 5 pixels 0-31 
assign ae_data_in_5b[5][0] = 5'b0;
assign ae_data_in_5b[5][1] = 5'b0;
assign ae_data_in_5b[5][2] = 5'b0;
assign ae_data_in_5b[5][3] = 5'b0;
assign ae_data_in_5b[5][4] = 5'b0;
assign ae_data_in_5b[5][5] = 5'b0;
assign ae_data_in_5b[5][6] = 5'b0;
assign ae_data_in_5b[5][7] = 5'b0;
assign ae_data_in_5b[5][8] = 5'b0;
assign ae_data_in_5b[5][9] = 5'b0;
assign ae_data_in_5b[5][10] = 5'b0;
assign ae_data_in_5b[5][11] = 5'b0;
assign ae_data_in_5b[5][12] = 5'b0;
assign ae_data_in_5b[5][13] = 5'b0;
assign ae_data_in_5b[5][14] = 5'b0;
assign ae_data_in_5b[5][15] = 5'b0;
assign ae_data_in_5b[5][16] = 5'b0;
assign ae_data_in_5b[5][17] = 5'b0;
assign ae_data_in_5b[5][18] = 5'b0;
assign ae_data_in_5b[5][19] = 5'b0;
assign ae_data_in_5b[5][20] = 5'b0;
assign ae_data_in_5b[5][21] = 5'b0;
assign ae_data_in_5b[5][22] = 5'b0;
assign ae_data_in_5b[5][23] = 5'b0;
assign ae_data_in_5b[5][24] = 5'b0;
assign ae_data_in_5b[5][25] = 5'b0;
assign ae_data_in_5b[5][26] = 5'b0;
assign ae_data_in_5b[5][27] = 5'b0;
assign ae_data_in_5b[5][28] = 5'b0;
assign ae_data_in_5b[5][29] = 5'b0;
assign ae_data_in_5b[5][30] = 5'b0;
assign ae_data_in_5b[5][31] = 5'b0;

// row 6 pixels 0-31 
assign ae_data_in_5b[6][0] = 5'b0;
assign ae_data_in_5b[6][1] = 5'b0;
assign ae_data_in_5b[6][2] = 5'b0;
assign ae_data_in_5b[6][3] = 5'b0;
assign ae_data_in_5b[6][4] = 5'b0;
assign ae_data_in_5b[6][5] = 5'b0;
assign ae_data_in_5b[6][6] = 5'b0;
assign ae_data_in_5b[6][7] = 5'b0;
assign ae_data_in_5b[6][8] = 5'b0;
assign ae_data_in_5b[6][9] = 5'b0;
assign ae_data_in_5b[6][10] = 5'b0;
assign ae_data_in_5b[6][11] = 5'b0;
assign ae_data_in_5b[6][12] = 5'b0;
assign ae_data_in_5b[6][13] = 5'b0;
assign ae_data_in_5b[6][14] = 5'b0;
assign ae_data_in_5b[6][15] = 5'b0;
assign ae_data_in_5b[6][16] = 5'b0;
assign ae_data_in_5b[6][17] = 5'b0;
assign ae_data_in_5b[6][18] = 5'b0;
assign ae_data_in_5b[6][19] = 5'b0;
assign ae_data_in_5b[6][20] = 5'b0;
assign ae_data_in_5b[6][21] = 5'b0;
assign ae_data_in_5b[6][22] = 5'b0;
assign ae_data_in_5b[6][23] = 5'b0;
assign ae_data_in_5b[6][24] = 5'b0;
assign ae_data_in_5b[6][25] = 5'b0;
assign ae_data_in_5b[6][26] = 5'b0;
assign ae_data_in_5b[6][27] = 5'b0;
assign ae_data_in_5b[6][28] = 5'b0;
assign ae_data_in_5b[6][29] = 5'b0;
assign ae_data_in_5b[6][30] = 5'b0;
assign ae_data_in_5b[6][31] = 5'b0;

// row 7 pixels 0-31 
assign ae_data_in_5b[7][0] = 5'b0;
assign ae_data_in_5b[7][1] = 5'b0;
assign ae_data_in_5b[7][2] = 5'b0;
assign ae_data_in_5b[7][3] = 5'b0;
assign ae_data_in_5b[7][4] = 5'b0;
assign ae_data_in_5b[7][5] = 5'b0;
assign ae_data_in_5b[7][6] = 5'b0;
assign ae_data_in_5b[7][7] = 5'b0;
assign ae_data_in_5b[7][8] = 5'b0;
assign ae_data_in_5b[7][9] = 5'b0;
assign ae_data_in_5b[7][10] = 5'b0;
assign ae_data_in_5b[7][11] = 5'b0;
assign ae_data_in_5b[7][12] = 5'b0;
assign ae_data_in_5b[7][13] = 5'b0;
assign ae_data_in_5b[7][14] = 5'b0;
assign ae_data_in_5b[7][15] = 5'b0;
assign ae_data_in_5b[7][16] = 5'b0;
assign ae_data_in_5b[7][17] = 5'b0;
assign ae_data_in_5b[7][18] = 5'b0;
assign ae_data_in_5b[7][19] = 5'b0;
assign ae_data_in_5b[7][20] = 5'b0;
assign ae_data_in_5b[7][21] = 5'b0;
assign ae_data_in_5b[7][22] = 5'b0;
assign ae_data_in_5b[7][23] = 5'b0;
assign ae_data_in_5b[7][24] = 5'b0;
assign ae_data_in_5b[7][25] = 5'b0;
assign ae_data_in_5b[7][26] = 5'b0;
assign ae_data_in_5b[7][27] = 5'b0;
assign ae_data_in_5b[7][28] = 5'b0;
assign ae_data_in_5b[7][29] = 5'b0;
assign ae_data_in_5b[7][30] = 5'b0;
assign ae_data_in_5b[7][31] = 5'b0;

// row 8 pixels 0-31 
assign ae_data_in_5b[8][0] = 5'b0;
assign ae_data_in_5b[8][1] = 5'b0;
assign ae_data_in_5b[8][2] = 5'b0;
assign ae_data_in_5b[8][3] = 5'b0;
assign ae_data_in_5b[8][4] = 5'b0;
assign ae_data_in_5b[8][5] = 5'b0;
assign ae_data_in_5b[8][6] = 5'b0;
assign ae_data_in_5b[8][7] = 5'b0;
assign ae_data_in_5b[8][8] = 5'b0;
assign ae_data_in_5b[8][9] = 5'b0;
assign ae_data_in_5b[8][10] = 5'b0;
assign ae_data_in_5b[8][11] = 5'b0;
assign ae_data_in_5b[8][12] = 5'b0;
assign ae_data_in_5b[8][13] = 5'b0;
assign ae_data_in_5b[8][14] = 5'b0;
assign ae_data_in_5b[8][15] = 5'b0;
assign ae_data_in_5b[8][16] = 5'b0;
assign ae_data_in_5b[8][17] = 5'b0;
assign ae_data_in_5b[8][18] = 5'b0;
assign ae_data_in_5b[8][19] = 5'b0;
assign ae_data_in_5b[8][20] = 5'b0;
assign ae_data_in_5b[8][21] = 5'b0;
assign ae_data_in_5b[8][22] = 5'b0;
assign ae_data_in_5b[8][23] = 5'b0;
assign ae_data_in_5b[8][24] = 5'b0;
assign ae_data_in_5b[8][25] = 5'b0;
assign ae_data_in_5b[8][26] = 5'b0;
assign ae_data_in_5b[8][27] = 5'b0;
assign ae_data_in_5b[8][28] = 5'b0;
assign ae_data_in_5b[8][29] = 5'b0;
assign ae_data_in_5b[8][30] = 5'b0;
assign ae_data_in_5b[8][31] = 5'b0;

// row 9 pixels 0-31 
assign ae_data_in_5b[9][0] = 5'b0;
assign ae_data_in_5b[9][1] = 5'b0;
assign ae_data_in_5b[9][2] = 5'b0;
assign ae_data_in_5b[9][3] = 5'b0;
assign ae_data_in_5b[9][4] = 5'b0;
assign ae_data_in_5b[9][5] = 5'b0;
assign ae_data_in_5b[9][6] = 5'b0;
assign ae_data_in_5b[9][7] = 5'b0;
assign ae_data_in_5b[9][8] = 5'b0;
assign ae_data_in_5b[9][9] = 5'b0;
assign ae_data_in_5b[9][10] = 5'b0;
assign ae_data_in_5b[9][11] = 5'b0;
assign ae_data_in_5b[9][12] = 5'b0;
assign ae_data_in_5b[9][13] = 5'b0;
assign ae_data_in_5b[9][14] = 5'b0;
assign ae_data_in_5b[9][15] = 5'b0;
assign ae_data_in_5b[9][16] = 5'b0;
assign ae_data_in_5b[9][17] = 5'b0;
assign ae_data_in_5b[9][18] = 5'b0;
assign ae_data_in_5b[9][19] = 5'b0;
assign ae_data_in_5b[9][20] = 5'b0;
assign ae_data_in_5b[9][21] = 5'b0;
assign ae_data_in_5b[9][22] = 5'b0;
assign ae_data_in_5b[9][23] = 5'b0;
assign ae_data_in_5b[9][24] = 5'b0;
assign ae_data_in_5b[9][25] = 5'b0;
assign ae_data_in_5b[9][26] = 5'b0;
assign ae_data_in_5b[9][27] = 5'b0;
assign ae_data_in_5b[9][28] = 5'b0;
assign ae_data_in_5b[9][29] = 5'b0;
assign ae_data_in_5b[9][30] = 5'b0;
assign ae_data_in_5b[9][31] = 5'b0;

// row 10 pixels 0-31 
assign ae_data_in_5b[10][0] = 5'b0;
assign ae_data_in_5b[10][1] = 5'b0;
assign ae_data_in_5b[10][2] = 5'b0;
assign ae_data_in_5b[10][3] = 5'b0;
assign ae_data_in_5b[10][4] = 5'b0;
assign ae_data_in_5b[10][5] = 5'b0;
assign ae_data_in_5b[10][6] = 5'b0;
assign ae_data_in_5b[10][7] = 5'b0;
assign ae_data_in_5b[10][8] = 5'b0;
assign ae_data_in_5b[10][9] = 5'b0;
assign ae_data_in_5b[10][10] = 5'b0;
assign ae_data_in_5b[10][11] = 5'b0;
assign ae_data_in_5b[10][12] = 5'b0;
assign ae_data_in_5b[10][13] = 5'b0;
assign ae_data_in_5b[10][14] = 5'b0;
assign ae_data_in_5b[10][15] = 5'b0;
assign ae_data_in_5b[10][16] = 5'b0;
assign ae_data_in_5b[10][17] = 5'b0;
assign ae_data_in_5b[10][18] = 5'b0;
assign ae_data_in_5b[10][19] = 5'b0;
assign ae_data_in_5b[10][20] = 5'b0;
assign ae_data_in_5b[10][21] = 5'b0;
assign ae_data_in_5b[10][22] = 5'b0;
assign ae_data_in_5b[10][23] = 5'b0;
assign ae_data_in_5b[10][24] = 5'b0;
assign ae_data_in_5b[10][25] = 5'b0;
assign ae_data_in_5b[10][26] = 5'b0;
assign ae_data_in_5b[10][27] = 5'b0;
assign ae_data_in_5b[10][28] = 5'b0;
assign ae_data_in_5b[10][29] = 5'b0;
assign ae_data_in_5b[10][30] = 5'b0;
assign ae_data_in_5b[10][31] = 5'b0;

// row 11 pixels 0-31 
assign ae_data_in_5b[11][0] = 5'b0;
assign ae_data_in_5b[11][1] = 5'b0;
assign ae_data_in_5b[11][2] = 5'b0;
assign ae_data_in_5b[11][3] = 5'b0;
assign ae_data_in_5b[11][4] = 5'b0;
assign ae_data_in_5b[11][5] = 5'b0;
assign ae_data_in_5b[11][6] = 5'b0;
assign ae_data_in_5b[11][7] = 5'b0;
assign ae_data_in_5b[11][8] = 5'b0;
assign ae_data_in_5b[11][9] = 5'b0;
assign ae_data_in_5b[11][10] = 5'b0;
assign ae_data_in_5b[11][11] = 5'b0;
assign ae_data_in_5b[11][12] = 5'b0;
assign ae_data_in_5b[11][13] = 5'b0;
assign ae_data_in_5b[11][14] = 5'b0;
assign ae_data_in_5b[11][15] = 5'b0;
assign ae_data_in_5b[11][16] = 5'b0;
assign ae_data_in_5b[11][17] = 5'b0;
assign ae_data_in_5b[11][18] = 5'b0;
assign ae_data_in_5b[11][19] = 5'b0;
assign ae_data_in_5b[11][20] = 5'b0;
assign ae_data_in_5b[11][21] = 5'b0;
assign ae_data_in_5b[11][22] = 5'b0;
assign ae_data_in_5b[11][23] = 5'b0;
assign ae_data_in_5b[11][24] = 5'b0;
assign ae_data_in_5b[11][25] = 5'b0;
assign ae_data_in_5b[11][26] = 5'b0;
assign ae_data_in_5b[11][27] = 5'b0;
assign ae_data_in_5b[11][28] = 5'b0;
assign ae_data_in_5b[11][29] = 5'b0;
assign ae_data_in_5b[11][30] = 5'b0;
assign ae_data_in_5b[11][31] = 5'b0;

// row 12 pixels 0-31 
assign ae_data_in_5b[12][0] = 5'b0;
assign ae_data_in_5b[12][1] = 5'b0;
assign ae_data_in_5b[12][2] = 5'b0;
assign ae_data_in_5b[12][3] = 5'b0;
assign ae_data_in_5b[12][4] = 5'b0;
assign ae_data_in_5b[12][5] = 5'b0;
assign ae_data_in_5b[12][6] = 5'b0;
assign ae_data_in_5b[12][7] = 5'b0;
assign ae_data_in_5b[12][8] = 5'b0;
assign ae_data_in_5b[12][9] = 5'b0;
assign ae_data_in_5b[12][10] = 5'b0;
assign ae_data_in_5b[12][11] = 5'b0;
assign ae_data_in_5b[12][12] = 5'b0;
assign ae_data_in_5b[12][13] = 5'b0;
assign ae_data_in_5b[12][14] = 5'b0;
assign ae_data_in_5b[12][15] = 5'b0;
assign ae_data_in_5b[12][16] = 5'b1;
assign ae_data_in_5b[12][17] = 5'b1;
assign ae_data_in_5b[12][18] = 5'b0;
assign ae_data_in_5b[12][19] = 5'b0;
assign ae_data_in_5b[12][20] = 5'b0;
assign ae_data_in_5b[12][21] = 5'b0;
assign ae_data_in_5b[12][22] = 5'b0;
assign ae_data_in_5b[12][23] = 5'b0;
assign ae_data_in_5b[12][24] = 5'b0;
assign ae_data_in_5b[12][25] = 5'b0;
assign ae_data_in_5b[12][26] = 5'b0;
assign ae_data_in_5b[12][27] = 5'b0;
assign ae_data_in_5b[12][28] = 5'b0;
assign ae_data_in_5b[12][29] = 5'b0;
assign ae_data_in_5b[12][30] = 5'b0;
assign ae_data_in_5b[12][31] = 5'b0;

// row 13 pixels 0-31 
assign ae_data_in_5b[13][0] = 5'b0;
assign ae_data_in_5b[13][1] = 5'b0;
assign ae_data_in_5b[13][2] = 5'b0;
assign ae_data_in_5b[13][3] = 5'b0;
assign ae_data_in_5b[13][4] = 5'b0;
assign ae_data_in_5b[13][5] = 5'b0;
assign ae_data_in_5b[13][6] = 5'b0;
assign ae_data_in_5b[13][7] = 5'b0;
assign ae_data_in_5b[13][8] = 5'b0;
assign ae_data_in_5b[13][9] = 5'b0;
assign ae_data_in_5b[13][10] = 5'b0;
assign ae_data_in_5b[13][11] = 5'b0;
assign ae_data_in_5b[13][12] = 5'b0;
assign ae_data_in_5b[13][13] = 5'b1;
assign ae_data_in_5b[13][14] = 5'b0;
assign ae_data_in_5b[13][15] = 5'b11;
assign ae_data_in_5b[13][16] = 5'b11;
assign ae_data_in_5b[13][17] = 5'b11;
assign ae_data_in_5b[13][18] = 5'b1;
assign ae_data_in_5b[13][19] = 5'b0;
assign ae_data_in_5b[13][20] = 5'b0;
assign ae_data_in_5b[13][21] = 5'b0;
assign ae_data_in_5b[13][22] = 5'b0;
assign ae_data_in_5b[13][23] = 5'b0;
assign ae_data_in_5b[13][24] = 5'b0;
assign ae_data_in_5b[13][25] = 5'b0;
assign ae_data_in_5b[13][26] = 5'b0;
assign ae_data_in_5b[13][27] = 5'b0;
assign ae_data_in_5b[13][28] = 5'b0;
assign ae_data_in_5b[13][29] = 5'b0;
assign ae_data_in_5b[13][30] = 5'b0;
assign ae_data_in_5b[13][31] = 5'b0;

// row 14 pixels 0-31 
assign ae_data_in_5b[14][0] = 5'b0;
assign ae_data_in_5b[14][1] = 5'b0;
assign ae_data_in_5b[14][2] = 5'b0;
assign ae_data_in_5b[14][3] = 5'b0;
assign ae_data_in_5b[14][4] = 5'b0;
assign ae_data_in_5b[14][5] = 5'b0;
assign ae_data_in_5b[14][6] = 5'b0;
assign ae_data_in_5b[14][7] = 5'b0;
assign ae_data_in_5b[14][8] = 5'b0;
assign ae_data_in_5b[14][9] = 5'b0;
assign ae_data_in_5b[14][10] = 5'b0;
assign ae_data_in_5b[14][11] = 5'b0;
assign ae_data_in_5b[14][12] = 5'b0;
assign ae_data_in_5b[14][13] = 5'b1;
assign ae_data_in_5b[14][14] = 5'b11;
assign ae_data_in_5b[14][15] = 5'b100;
assign ae_data_in_5b[14][16] = 5'b1000;
assign ae_data_in_5b[14][17] = 5'b101;
assign ae_data_in_5b[14][18] = 5'b11;
assign ae_data_in_5b[14][19] = 5'b0;
assign ae_data_in_5b[14][20] = 5'b0;
assign ae_data_in_5b[14][21] = 5'b0;
assign ae_data_in_5b[14][22] = 5'b0;
assign ae_data_in_5b[14][23] = 5'b0;
assign ae_data_in_5b[14][24] = 5'b0;
assign ae_data_in_5b[14][25] = 5'b0;
assign ae_data_in_5b[14][26] = 5'b0;
assign ae_data_in_5b[14][27] = 5'b0;
assign ae_data_in_5b[14][28] = 5'b0;
assign ae_data_in_5b[14][29] = 5'b0;
assign ae_data_in_5b[14][30] = 5'b0;
assign ae_data_in_5b[14][31] = 5'b0;

// row 15 pixels 0-31 
assign ae_data_in_5b[15][0] = 5'b0;
assign ae_data_in_5b[15][1] = 5'b0;
assign ae_data_in_5b[15][2] = 5'b0;
assign ae_data_in_5b[15][3] = 5'b0;
assign ae_data_in_5b[15][4] = 5'b0;
assign ae_data_in_5b[15][5] = 5'b0;
assign ae_data_in_5b[15][6] = 5'b0;
assign ae_data_in_5b[15][7] = 5'b0;
assign ae_data_in_5b[15][8] = 5'b0;
assign ae_data_in_5b[15][9] = 5'b0;
assign ae_data_in_5b[15][10] = 5'b0;
assign ae_data_in_5b[15][11] = 5'b0;
assign ae_data_in_5b[15][12] = 5'b0;
assign ae_data_in_5b[15][13] = 5'b1;
assign ae_data_in_5b[15][14] = 5'b101;
assign ae_data_in_5b[15][15] = 5'b10001;
assign ae_data_in_5b[15][16] = 5'b10110;
assign ae_data_in_5b[15][17] = 5'b10011;
assign ae_data_in_5b[15][18] = 5'b101;
assign ae_data_in_5b[15][19] = 5'b11;
assign ae_data_in_5b[15][20] = 5'b0;
assign ae_data_in_5b[15][21] = 5'b0;
assign ae_data_in_5b[15][22] = 5'b0;
assign ae_data_in_5b[15][23] = 5'b0;
assign ae_data_in_5b[15][24] = 5'b0;
assign ae_data_in_5b[15][25] = 5'b0;
assign ae_data_in_5b[15][26] = 5'b0;
assign ae_data_in_5b[15][27] = 5'b0;
assign ae_data_in_5b[15][28] = 5'b0;
assign ae_data_in_5b[15][29] = 5'b0;
assign ae_data_in_5b[15][30] = 5'b0;
assign ae_data_in_5b[15][31] = 5'b0;

// row 16 pixels 0-31 
assign ae_data_in_5b[16][0] = 5'b0;
assign ae_data_in_5b[16][1] = 5'b0;
assign ae_data_in_5b[16][2] = 5'b0;
assign ae_data_in_5b[16][3] = 5'b0;
assign ae_data_in_5b[16][4] = 5'b0;
assign ae_data_in_5b[16][5] = 5'b0;
assign ae_data_in_5b[16][6] = 5'b0;
assign ae_data_in_5b[16][7] = 5'b0;
assign ae_data_in_5b[16][8] = 5'b0;
assign ae_data_in_5b[16][9] = 5'b0;
assign ae_data_in_5b[16][10] = 5'b0;
assign ae_data_in_5b[16][11] = 5'b0;
assign ae_data_in_5b[16][12] = 5'b1;
assign ae_data_in_5b[16][13] = 5'b11;
assign ae_data_in_5b[16][14] = 5'b1000;
assign ae_data_in_5b[16][15] = 5'b10110;
assign ae_data_in_5b[16][16] = 5'b11100;
assign ae_data_in_5b[16][17] = 5'b10110;
assign ae_data_in_5b[16][18] = 5'b1000;
assign ae_data_in_5b[16][19] = 5'b11;
assign ae_data_in_5b[16][20] = 5'b0;
assign ae_data_in_5b[16][21] = 5'b0;
assign ae_data_in_5b[16][22] = 5'b0;
assign ae_data_in_5b[16][23] = 5'b0;
assign ae_data_in_5b[16][24] = 5'b0;
assign ae_data_in_5b[16][25] = 5'b0;
assign ae_data_in_5b[16][26] = 5'b0;
assign ae_data_in_5b[16][27] = 5'b0;
assign ae_data_in_5b[16][28] = 5'b0;
assign ae_data_in_5b[16][29] = 5'b0;
assign ae_data_in_5b[16][30] = 5'b0;
assign ae_data_in_5b[16][31] = 5'b0;

// row 17 pixels 0-31 
assign ae_data_in_5b[17][0] = 5'b0;
assign ae_data_in_5b[17][1] = 5'b0;
assign ae_data_in_5b[17][2] = 5'b0;
assign ae_data_in_5b[17][3] = 5'b0;
assign ae_data_in_5b[17][4] = 5'b0;
assign ae_data_in_5b[17][5] = 5'b0;
assign ae_data_in_5b[17][6] = 5'b0;
assign ae_data_in_5b[17][7] = 5'b0;
assign ae_data_in_5b[17][8] = 5'b0;
assign ae_data_in_5b[17][9] = 5'b0;
assign ae_data_in_5b[17][10] = 5'b0;
assign ae_data_in_5b[17][11] = 5'b0;
assign ae_data_in_5b[17][12] = 5'b0;
assign ae_data_in_5b[17][13] = 5'b10;
assign ae_data_in_5b[17][14] = 5'b101;
assign ae_data_in_5b[17][15] = 5'b10010;
assign ae_data_in_5b[17][16] = 5'b10110;
assign ae_data_in_5b[17][17] = 5'b10010;
assign ae_data_in_5b[17][18] = 5'b101;
assign ae_data_in_5b[17][19] = 5'b10;
assign ae_data_in_5b[17][20] = 5'b0;
assign ae_data_in_5b[17][21] = 5'b0;
assign ae_data_in_5b[17][22] = 5'b0;
assign ae_data_in_5b[17][23] = 5'b0;
assign ae_data_in_5b[17][24] = 5'b0;
assign ae_data_in_5b[17][25] = 5'b0;
assign ae_data_in_5b[17][26] = 5'b0;
assign ae_data_in_5b[17][27] = 5'b0;
assign ae_data_in_5b[17][28] = 5'b0;
assign ae_data_in_5b[17][29] = 5'b0;
assign ae_data_in_5b[17][30] = 5'b0;
assign ae_data_in_5b[17][31] = 5'b0;

// row 18 pixels 0-31 
assign ae_data_in_5b[18][0] = 5'b0;
assign ae_data_in_5b[18][1] = 5'b0;
assign ae_data_in_5b[18][2] = 5'b0;
assign ae_data_in_5b[18][3] = 5'b0;
assign ae_data_in_5b[18][4] = 5'b0;
assign ae_data_in_5b[18][5] = 5'b0;
assign ae_data_in_5b[18][6] = 5'b0;
assign ae_data_in_5b[18][7] = 5'b0;
assign ae_data_in_5b[18][8] = 5'b0;
assign ae_data_in_5b[18][9] = 5'b0;
assign ae_data_in_5b[18][10] = 5'b0;
assign ae_data_in_5b[18][11] = 5'b0;
assign ae_data_in_5b[18][12] = 5'b0;
assign ae_data_in_5b[18][13] = 5'b10;
assign ae_data_in_5b[18][14] = 5'b11;
assign ae_data_in_5b[18][15] = 5'b101;
assign ae_data_in_5b[18][16] = 5'b1000;
assign ae_data_in_5b[18][17] = 5'b101;
assign ae_data_in_5b[18][18] = 5'b11;
assign ae_data_in_5b[18][19] = 5'b1;
assign ae_data_in_5b[18][20] = 5'b0;
assign ae_data_in_5b[18][21] = 5'b0;
assign ae_data_in_5b[18][22] = 5'b0;
assign ae_data_in_5b[18][23] = 5'b0;
assign ae_data_in_5b[18][24] = 5'b0;
assign ae_data_in_5b[18][25] = 5'b0;
assign ae_data_in_5b[18][26] = 5'b0;
assign ae_data_in_5b[18][27] = 5'b0;
assign ae_data_in_5b[18][28] = 5'b0;
assign ae_data_in_5b[18][29] = 5'b0;
assign ae_data_in_5b[18][30] = 5'b0;
assign ae_data_in_5b[18][31] = 5'b0;

// row 19 pixels 0-31 
assign ae_data_in_5b[19][0] = 5'b0;
assign ae_data_in_5b[19][1] = 5'b0;
assign ae_data_in_5b[19][2] = 5'b0;
assign ae_data_in_5b[19][3] = 5'b0;
assign ae_data_in_5b[19][4] = 5'b0;
assign ae_data_in_5b[19][5] = 5'b0;
assign ae_data_in_5b[19][6] = 5'b0;
assign ae_data_in_5b[19][7] = 5'b0;
assign ae_data_in_5b[19][8] = 5'b0;
assign ae_data_in_5b[19][9] = 5'b0;
assign ae_data_in_5b[19][10] = 5'b0;
assign ae_data_in_5b[19][11] = 5'b0;
assign ae_data_in_5b[19][12] = 5'b0;
assign ae_data_in_5b[19][13] = 5'b0;
assign ae_data_in_5b[19][14] = 5'b0;
assign ae_data_in_5b[19][15] = 5'b11;
assign ae_data_in_5b[19][16] = 5'b11;
assign ae_data_in_5b[19][17] = 5'b10;
assign ae_data_in_5b[19][18] = 5'b0;
assign ae_data_in_5b[19][19] = 5'b0;
assign ae_data_in_5b[19][20] = 5'b0;
assign ae_data_in_5b[19][21] = 5'b0;
assign ae_data_in_5b[19][22] = 5'b0;
assign ae_data_in_5b[19][23] = 5'b0;
assign ae_data_in_5b[19][24] = 5'b0;
assign ae_data_in_5b[19][25] = 5'b0;
assign ae_data_in_5b[19][26] = 5'b0;
assign ae_data_in_5b[19][27] = 5'b0;
assign ae_data_in_5b[19][28] = 5'b0;
assign ae_data_in_5b[19][29] = 5'b0;
assign ae_data_in_5b[19][30] = 5'b0;
assign ae_data_in_5b[19][31] = 5'b0;

// row 20 pixels 0-31 
assign ae_data_in_5b[20][0] = 5'b0;
assign ae_data_in_5b[20][1] = 5'b0;
assign ae_data_in_5b[20][2] = 5'b0;
assign ae_data_in_5b[20][3] = 5'b0;
assign ae_data_in_5b[20][4] = 5'b0;
assign ae_data_in_5b[20][5] = 5'b0;
assign ae_data_in_5b[20][6] = 5'b0;
assign ae_data_in_5b[20][7] = 5'b0;
assign ae_data_in_5b[20][8] = 5'b0;
assign ae_data_in_5b[20][9] = 5'b0;
assign ae_data_in_5b[20][10] = 5'b0;
assign ae_data_in_5b[20][11] = 5'b0;
assign ae_data_in_5b[20][12] = 5'b0;
assign ae_data_in_5b[20][13] = 5'b0;
assign ae_data_in_5b[20][14] = 5'b1;
assign ae_data_in_5b[20][15] = 5'b0;
assign ae_data_in_5b[20][16] = 5'b1;
assign ae_data_in_5b[20][17] = 5'b0;
assign ae_data_in_5b[20][18] = 5'b0;
assign ae_data_in_5b[20][19] = 5'b0;
assign ae_data_in_5b[20][20] = 5'b0;
assign ae_data_in_5b[20][21] = 5'b0;
assign ae_data_in_5b[20][22] = 5'b0;
assign ae_data_in_5b[20][23] = 5'b0;
assign ae_data_in_5b[20][24] = 5'b0;
assign ae_data_in_5b[20][25] = 5'b0;
assign ae_data_in_5b[20][26] = 5'b0;
assign ae_data_in_5b[20][27] = 5'b0;
assign ae_data_in_5b[20][28] = 5'b0;
assign ae_data_in_5b[20][29] = 5'b0;
assign ae_data_in_5b[20][30] = 5'b0;
assign ae_data_in_5b[20][31] = 5'b0;

// row 21 pixels 0-31 
assign ae_data_in_5b[21][0] = 5'b0;
assign ae_data_in_5b[21][1] = 5'b0;
assign ae_data_in_5b[21][2] = 5'b0;
assign ae_data_in_5b[21][3] = 5'b0;
assign ae_data_in_5b[21][4] = 5'b0;
assign ae_data_in_5b[21][5] = 5'b0;
assign ae_data_in_5b[21][6] = 5'b0;
assign ae_data_in_5b[21][7] = 5'b0;
assign ae_data_in_5b[21][8] = 5'b0;
assign ae_data_in_5b[21][9] = 5'b0;
assign ae_data_in_5b[21][10] = 5'b0;
assign ae_data_in_5b[21][11] = 5'b0;
assign ae_data_in_5b[21][12] = 5'b0;
assign ae_data_in_5b[21][13] = 5'b0;
assign ae_data_in_5b[21][14] = 5'b0;
assign ae_data_in_5b[21][15] = 5'b1;
assign ae_data_in_5b[21][16] = 5'b0;
assign ae_data_in_5b[21][17] = 5'b0;
assign ae_data_in_5b[21][18] = 5'b0;
assign ae_data_in_5b[21][19] = 5'b0;
assign ae_data_in_5b[21][20] = 5'b0;
assign ae_data_in_5b[21][21] = 5'b0;
assign ae_data_in_5b[21][22] = 5'b0;
assign ae_data_in_5b[21][23] = 5'b0;
assign ae_data_in_5b[21][24] = 5'b0;
assign ae_data_in_5b[21][25] = 5'b0;
assign ae_data_in_5b[21][26] = 5'b0;
assign ae_data_in_5b[21][27] = 5'b0;
assign ae_data_in_5b[21][28] = 5'b0;
assign ae_data_in_5b[21][29] = 5'b0;
assign ae_data_in_5b[21][30] = 5'b0;
assign ae_data_in_5b[21][31] = 5'b0;

// row 22 pixels 0-31 
assign ae_data_in_5b[22][0] = 5'b0;
assign ae_data_in_5b[22][1] = 5'b0;
assign ae_data_in_5b[22][2] = 5'b0;
assign ae_data_in_5b[22][3] = 5'b0;
assign ae_data_in_5b[22][4] = 5'b0;
assign ae_data_in_5b[22][5] = 5'b0;
assign ae_data_in_5b[22][6] = 5'b0;
assign ae_data_in_5b[22][7] = 5'b0;
assign ae_data_in_5b[22][8] = 5'b0;
assign ae_data_in_5b[22][9] = 5'b0;
assign ae_data_in_5b[22][10] = 5'b0;
assign ae_data_in_5b[22][11] = 5'b0;
assign ae_data_in_5b[22][12] = 5'b0;
assign ae_data_in_5b[22][13] = 5'b0;
assign ae_data_in_5b[22][14] = 5'b0;
assign ae_data_in_5b[22][15] = 5'b0;
assign ae_data_in_5b[22][16] = 5'b0;
assign ae_data_in_5b[22][17] = 5'b0;
assign ae_data_in_5b[22][18] = 5'b0;
assign ae_data_in_5b[22][19] = 5'b0;
assign ae_data_in_5b[22][20] = 5'b0;
assign ae_data_in_5b[22][21] = 5'b0;
assign ae_data_in_5b[22][22] = 5'b0;
assign ae_data_in_5b[22][23] = 5'b0;
assign ae_data_in_5b[22][24] = 5'b0;
assign ae_data_in_5b[22][25] = 5'b0;
assign ae_data_in_5b[22][26] = 5'b0;
assign ae_data_in_5b[22][27] = 5'b0;
assign ae_data_in_5b[22][28] = 5'b0;
assign ae_data_in_5b[22][29] = 5'b0;
assign ae_data_in_5b[22][30] = 5'b0;
assign ae_data_in_5b[22][31] = 5'b0;

// row 23 pixels 0-31 
assign ae_data_in_5b[23][0] = 5'b0;
assign ae_data_in_5b[23][1] = 5'b0;
assign ae_data_in_5b[23][2] = 5'b0;
assign ae_data_in_5b[23][3] = 5'b0;
assign ae_data_in_5b[23][4] = 5'b0;
assign ae_data_in_5b[23][5] = 5'b0;
assign ae_data_in_5b[23][6] = 5'b0;
assign ae_data_in_5b[23][7] = 5'b0;
assign ae_data_in_5b[23][8] = 5'b0;
assign ae_data_in_5b[23][9] = 5'b0;
assign ae_data_in_5b[23][10] = 5'b0;
assign ae_data_in_5b[23][11] = 5'b0;
assign ae_data_in_5b[23][12] = 5'b0;
assign ae_data_in_5b[23][13] = 5'b0;
assign ae_data_in_5b[23][14] = 5'b0;
assign ae_data_in_5b[23][15] = 5'b0;
assign ae_data_in_5b[23][16] = 5'b0;
assign ae_data_in_5b[23][17] = 5'b0;
assign ae_data_in_5b[23][18] = 5'b0;
assign ae_data_in_5b[23][19] = 5'b0;
assign ae_data_in_5b[23][20] = 5'b0;
assign ae_data_in_5b[23][21] = 5'b0;
assign ae_data_in_5b[23][22] = 5'b0;
assign ae_data_in_5b[23][23] = 5'b0;
assign ae_data_in_5b[23][24] = 5'b0;
assign ae_data_in_5b[23][25] = 5'b0;
assign ae_data_in_5b[23][26] = 5'b0;
assign ae_data_in_5b[23][27] = 5'b0;
assign ae_data_in_5b[23][28] = 5'b0;
assign ae_data_in_5b[23][29] = 5'b0;
assign ae_data_in_5b[23][30] = 5'b0;
assign ae_data_in_5b[23][31] = 5'b0;

// row 24 pixels 0-31 
assign ae_data_in_5b[24][0] = 5'b0;
assign ae_data_in_5b[24][1] = 5'b0;
assign ae_data_in_5b[24][2] = 5'b0;
assign ae_data_in_5b[24][3] = 5'b0;
assign ae_data_in_5b[24][4] = 5'b0;
assign ae_data_in_5b[24][5] = 5'b0;
assign ae_data_in_5b[24][6] = 5'b0;
assign ae_data_in_5b[24][7] = 5'b0;
assign ae_data_in_5b[24][8] = 5'b0;
assign ae_data_in_5b[24][9] = 5'b0;
assign ae_data_in_5b[24][10] = 5'b0;
assign ae_data_in_5b[24][11] = 5'b0;
assign ae_data_in_5b[24][12] = 5'b0;
assign ae_data_in_5b[24][13] = 5'b0;
assign ae_data_in_5b[24][14] = 5'b0;
assign ae_data_in_5b[24][15] = 5'b0;
assign ae_data_in_5b[24][16] = 5'b0;
assign ae_data_in_5b[24][17] = 5'b0;
assign ae_data_in_5b[24][18] = 5'b0;
assign ae_data_in_5b[24][19] = 5'b0;
assign ae_data_in_5b[24][20] = 5'b0;
assign ae_data_in_5b[24][21] = 5'b0;
assign ae_data_in_5b[24][22] = 5'b0;
assign ae_data_in_5b[24][23] = 5'b0;
assign ae_data_in_5b[24][24] = 5'b0;
assign ae_data_in_5b[24][25] = 5'b0;
assign ae_data_in_5b[24][26] = 5'b0;
assign ae_data_in_5b[24][27] = 5'b0;
assign ae_data_in_5b[24][28] = 5'b0;
assign ae_data_in_5b[24][29] = 5'b0;
assign ae_data_in_5b[24][30] = 5'b0;
assign ae_data_in_5b[24][31] = 5'b0;

// row 25 pixels 0-31 
assign ae_data_in_5b[25][0] = 5'b0;
assign ae_data_in_5b[25][1] = 5'b0;
assign ae_data_in_5b[25][2] = 5'b0;
assign ae_data_in_5b[25][3] = 5'b0;
assign ae_data_in_5b[25][4] = 5'b0;
assign ae_data_in_5b[25][5] = 5'b0;
assign ae_data_in_5b[25][6] = 5'b0;
assign ae_data_in_5b[25][7] = 5'b0;
assign ae_data_in_5b[25][8] = 5'b0;
assign ae_data_in_5b[25][9] = 5'b0;
assign ae_data_in_5b[25][10] = 5'b0;
assign ae_data_in_5b[25][11] = 5'b0;
assign ae_data_in_5b[25][12] = 5'b0;
assign ae_data_in_5b[25][13] = 5'b0;
assign ae_data_in_5b[25][14] = 5'b0;
assign ae_data_in_5b[25][15] = 5'b0;
assign ae_data_in_5b[25][16] = 5'b0;
assign ae_data_in_5b[25][17] = 5'b0;
assign ae_data_in_5b[25][18] = 5'b0;
assign ae_data_in_5b[25][19] = 5'b0;
assign ae_data_in_5b[25][20] = 5'b0;
assign ae_data_in_5b[25][21] = 5'b0;
assign ae_data_in_5b[25][22] = 5'b0;
assign ae_data_in_5b[25][23] = 5'b0;
assign ae_data_in_5b[25][24] = 5'b0;
assign ae_data_in_5b[25][25] = 5'b0;
assign ae_data_in_5b[25][26] = 5'b0;
assign ae_data_in_5b[25][27] = 5'b0;
assign ae_data_in_5b[25][28] = 5'b0;
assign ae_data_in_5b[25][29] = 5'b0;
assign ae_data_in_5b[25][30] = 5'b0;
assign ae_data_in_5b[25][31] = 5'b0;

// row 26 pixels 0-31 
assign ae_data_in_5b[26][0] = 5'b0;
assign ae_data_in_5b[26][1] = 5'b0;
assign ae_data_in_5b[26][2] = 5'b0;
assign ae_data_in_5b[26][3] = 5'b0;
assign ae_data_in_5b[26][4] = 5'b0;
assign ae_data_in_5b[26][5] = 5'b0;
assign ae_data_in_5b[26][6] = 5'b0;
assign ae_data_in_5b[26][7] = 5'b0;
assign ae_data_in_5b[26][8] = 5'b0;
assign ae_data_in_5b[26][9] = 5'b0;
assign ae_data_in_5b[26][10] = 5'b0;
assign ae_data_in_5b[26][11] = 5'b0;
assign ae_data_in_5b[26][12] = 5'b0;
assign ae_data_in_5b[26][13] = 5'b0;
assign ae_data_in_5b[26][14] = 5'b0;
assign ae_data_in_5b[26][15] = 5'b0;
assign ae_data_in_5b[26][16] = 5'b0;
assign ae_data_in_5b[26][17] = 5'b0;
assign ae_data_in_5b[26][18] = 5'b0;
assign ae_data_in_5b[26][19] = 5'b0;
assign ae_data_in_5b[26][20] = 5'b0;
assign ae_data_in_5b[26][21] = 5'b0;
assign ae_data_in_5b[26][22] = 5'b0;
assign ae_data_in_5b[26][23] = 5'b0;
assign ae_data_in_5b[26][24] = 5'b0;
assign ae_data_in_5b[26][25] = 5'b0;
assign ae_data_in_5b[26][26] = 5'b0;
assign ae_data_in_5b[26][27] = 5'b0;
assign ae_data_in_5b[26][28] = 5'b0;
assign ae_data_in_5b[26][29] = 5'b0;
assign ae_data_in_5b[26][30] = 5'b0;
assign ae_data_in_5b[26][31] = 5'b0;

// row 27 pixels 0-31 
assign ae_data_in_5b[27][0] = 5'b0;
assign ae_data_in_5b[27][1] = 5'b0;
assign ae_data_in_5b[27][2] = 5'b0;
assign ae_data_in_5b[27][3] = 5'b0;
assign ae_data_in_5b[27][4] = 5'b0;
assign ae_data_in_5b[27][5] = 5'b0;
assign ae_data_in_5b[27][6] = 5'b0;
assign ae_data_in_5b[27][7] = 5'b0;
assign ae_data_in_5b[27][8] = 5'b0;
assign ae_data_in_5b[27][9] = 5'b0;
assign ae_data_in_5b[27][10] = 5'b0;
assign ae_data_in_5b[27][11] = 5'b0;
assign ae_data_in_5b[27][12] = 5'b0;
assign ae_data_in_5b[27][13] = 5'b0;
assign ae_data_in_5b[27][14] = 5'b0;
assign ae_data_in_5b[27][15] = 5'b0;
assign ae_data_in_5b[27][16] = 5'b0;
assign ae_data_in_5b[27][17] = 5'b0;
assign ae_data_in_5b[27][18] = 5'b0;
assign ae_data_in_5b[27][19] = 5'b0;
assign ae_data_in_5b[27][20] = 5'b0;
assign ae_data_in_5b[27][21] = 5'b0;
assign ae_data_in_5b[27][22] = 5'b0;
assign ae_data_in_5b[27][23] = 5'b0;
assign ae_data_in_5b[27][24] = 5'b0;
assign ae_data_in_5b[27][25] = 5'b0;
assign ae_data_in_5b[27][26] = 5'b0;
assign ae_data_in_5b[27][27] = 5'b0;
assign ae_data_in_5b[27][28] = 5'b0;
assign ae_data_in_5b[27][29] = 5'b0;
assign ae_data_in_5b[27][30] = 5'b0;
assign ae_data_in_5b[27][31] = 5'b0;

// row 28 pixels 0-31 
assign ae_data_in_5b[28][0] = 5'b0;
assign ae_data_in_5b[28][1] = 5'b0;
assign ae_data_in_5b[28][2] = 5'b0;
assign ae_data_in_5b[28][3] = 5'b0;
assign ae_data_in_5b[28][4] = 5'b0;
assign ae_data_in_5b[28][5] = 5'b0;
assign ae_data_in_5b[28][6] = 5'b0;
assign ae_data_in_5b[28][7] = 5'b0;
assign ae_data_in_5b[28][8] = 5'b0;
assign ae_data_in_5b[28][9] = 5'b0;
assign ae_data_in_5b[28][10] = 5'b0;
assign ae_data_in_5b[28][11] = 5'b0;
assign ae_data_in_5b[28][12] = 5'b0;
assign ae_data_in_5b[28][13] = 5'b0;
assign ae_data_in_5b[28][14] = 5'b0;
assign ae_data_in_5b[28][15] = 5'b0;
assign ae_data_in_5b[28][16] = 5'b0;
assign ae_data_in_5b[28][17] = 5'b0;
assign ae_data_in_5b[28][18] = 5'b0;
assign ae_data_in_5b[28][19] = 5'b0;
assign ae_data_in_5b[28][20] = 5'b0;
assign ae_data_in_5b[28][21] = 5'b0;
assign ae_data_in_5b[28][22] = 5'b0;
assign ae_data_in_5b[28][23] = 5'b0;
assign ae_data_in_5b[28][24] = 5'b0;
assign ae_data_in_5b[28][25] = 5'b0;
assign ae_data_in_5b[28][26] = 5'b0;
assign ae_data_in_5b[28][27] = 5'b0;
assign ae_data_in_5b[28][28] = 5'b0;
assign ae_data_in_5b[28][29] = 5'b0;
assign ae_data_in_5b[28][30] = 5'b0;
assign ae_data_in_5b[28][31] = 5'b0;

// row 29 pixels 0-31 
assign ae_data_in_5b[29][0] = 5'b0;
assign ae_data_in_5b[29][1] = 5'b0;
assign ae_data_in_5b[29][2] = 5'b0;
assign ae_data_in_5b[29][3] = 5'b0;
assign ae_data_in_5b[29][4] = 5'b0;
assign ae_data_in_5b[29][5] = 5'b0;
assign ae_data_in_5b[29][6] = 5'b0;
assign ae_data_in_5b[29][7] = 5'b0;
assign ae_data_in_5b[29][8] = 5'b0;
assign ae_data_in_5b[29][9] = 5'b0;
assign ae_data_in_5b[29][10] = 5'b0;
assign ae_data_in_5b[29][11] = 5'b0;
assign ae_data_in_5b[29][12] = 5'b0;
assign ae_data_in_5b[29][13] = 5'b0;
assign ae_data_in_5b[29][14] = 5'b0;
assign ae_data_in_5b[29][15] = 5'b0;
assign ae_data_in_5b[29][16] = 5'b0;
assign ae_data_in_5b[29][17] = 5'b0;
assign ae_data_in_5b[29][18] = 5'b0;
assign ae_data_in_5b[29][19] = 5'b0;
assign ae_data_in_5b[29][20] = 5'b0;
assign ae_data_in_5b[29][21] = 5'b0;
assign ae_data_in_5b[29][22] = 5'b0;
assign ae_data_in_5b[29][23] = 5'b0;
assign ae_data_in_5b[29][24] = 5'b0;
assign ae_data_in_5b[29][25] = 5'b0;
assign ae_data_in_5b[29][26] = 5'b0;
assign ae_data_in_5b[29][27] = 5'b0;
assign ae_data_in_5b[29][28] = 5'b0;
assign ae_data_in_5b[29][29] = 5'b0;
assign ae_data_in_5b[29][30] = 5'b0;
assign ae_data_in_5b[29][31] = 5'b0;

// row 30 pixels 0-31 
assign ae_data_in_5b[30][0] = 5'b0;
assign ae_data_in_5b[30][1] = 5'b0;
assign ae_data_in_5b[30][2] = 5'b0;
assign ae_data_in_5b[30][3] = 5'b0;
assign ae_data_in_5b[30][4] = 5'b0;
assign ae_data_in_5b[30][5] = 5'b0;
assign ae_data_in_5b[30][6] = 5'b0;
assign ae_data_in_5b[30][7] = 5'b0;
assign ae_data_in_5b[30][8] = 5'b0;
assign ae_data_in_5b[30][9] = 5'b0;
assign ae_data_in_5b[30][10] = 5'b0;
assign ae_data_in_5b[30][11] = 5'b0;
assign ae_data_in_5b[30][12] = 5'b0;
assign ae_data_in_5b[30][13] = 5'b0;
assign ae_data_in_5b[30][14] = 5'b0;
assign ae_data_in_5b[30][15] = 5'b0;
assign ae_data_in_5b[30][16] = 5'b0;
assign ae_data_in_5b[30][17] = 5'b0;
assign ae_data_in_5b[30][18] = 5'b0;
assign ae_data_in_5b[30][19] = 5'b0;
assign ae_data_in_5b[30][20] = 5'b0;
assign ae_data_in_5b[30][21] = 5'b0;
assign ae_data_in_5b[30][22] = 5'b0;
assign ae_data_in_5b[30][23] = 5'b0;
assign ae_data_in_5b[30][24] = 5'b0;
assign ae_data_in_5b[30][25] = 5'b0;
assign ae_data_in_5b[30][26] = 5'b0;
assign ae_data_in_5b[30][27] = 5'b0;
assign ae_data_in_5b[30][28] = 5'b0;
assign ae_data_in_5b[30][29] = 5'b0;
assign ae_data_in_5b[30][30] = 5'b0;
assign ae_data_in_5b[30][31] = 5'b0;

// row 31 pixels 0-31 
assign ae_data_in_5b[31][0] = 5'b0;
assign ae_data_in_5b[31][1] = 5'b0;
assign ae_data_in_5b[31][2] = 5'b0;
assign ae_data_in_5b[31][3] = 5'b0;
assign ae_data_in_5b[31][4] = 5'b0;
assign ae_data_in_5b[31][5] = 5'b0;
assign ae_data_in_5b[31][6] = 5'b0;
assign ae_data_in_5b[31][7] = 5'b0;
assign ae_data_in_5b[31][8] = 5'b0;
assign ae_data_in_5b[31][9] = 5'b0;
assign ae_data_in_5b[31][10] = 5'b0;
assign ae_data_in_5b[31][11] = 5'b0;
assign ae_data_in_5b[31][12] = 5'b0;
assign ae_data_in_5b[31][13] = 5'b0;
assign ae_data_in_5b[31][14] = 5'b0;
assign ae_data_in_5b[31][15] = 5'b0;
assign ae_data_in_5b[31][16] = 5'b0;
assign ae_data_in_5b[31][17] = 5'b0;
assign ae_data_in_5b[31][18] = 5'b0;
assign ae_data_in_5b[31][19] = 5'b0;
assign ae_data_in_5b[31][20] = 5'b0;
assign ae_data_in_5b[31][21] = 5'b0;
assign ae_data_in_5b[31][22] = 5'b0;
assign ae_data_in_5b[31][23] = 5'b0;
assign ae_data_in_5b[31][24] = 5'b0;
assign ae_data_in_5b[31][25] = 5'b0;
assign ae_data_in_5b[31][26] = 5'b0;
assign ae_data_in_5b[31][27] = 5'b0;
assign ae_data_in_5b[31][28] = 5'b0;
assign ae_data_in_5b[31][29] = 5'b0;
assign ae_data_in_5b[31][30] = 5'b0;
assign ae_data_in_5b[31][31] = 5'b0;



// 19b PCA outputs 

assign pca_output_19b[0] = 19'b1100010101000100001;
assign pca_output_19b[1] = 19'b1111111110111111111;
assign pca_output_19b[2] = 19'b11011100001;
assign pca_output_19b[3] = 19'b1111111110101010101;
assign pca_output_19b[4] = 19'b1111111111011000111;
assign pca_output_19b[5] = 19'b1111111101010100000;
assign pca_output_19b[6] = 19'b1111111111110111111;
assign pca_output_19b[7] = 19'b111011101;
assign pca_output_19b[8] = 19'b1010010000;
assign pca_output_19b[9] = 19'b1111111110000011101;
assign pca_output_19b[10] = 19'b1011101;
assign pca_output_19b[11] = 19'b1111111111000100100;
assign pca_output_19b[12] = 19'b1000111010;
assign pca_output_19b[13] = 19'b1010101111;
assign pca_output_19b[14] = 19'b1111111011101100010;
assign pca_output_19b[15] = 19'b101010101;
assign pca_output_19b[16] = 19'b1111111110011001011;
assign pca_output_19b[17] = 19'b11101110110;
assign pca_output_19b[18] = 19'b1111111110111010001;
assign pca_output_19b[19] = 19'b10110110;
assign pca_output_19b[20] = 19'b1111111110110110000;
assign pca_output_19b[21] = 19'b1111111111101010110;
assign pca_output_19b[22] = 19'b1111111111011010001;
assign pca_output_19b[23] = 19'b111;
assign pca_output_19b[24] = 19'b1010;
assign pca_output_19b[25] = 19'b1000000;
assign pca_output_19b[26] = 19'b1111111111110111010;
assign pca_output_19b[27] = 19'b111101111;
assign pca_output_19b[28] = 19'b1111111111001000100;
assign pca_output_19b[29] = 19'b1111111111110111000;



// 5b AE outputs 

assign ae_output_5b[0] = 5'b0;
assign ae_output_5b[1] = 5'b11110;
assign ae_output_5b[2] = 5'b11010;
assign ae_output_5b[3] = 5'b11111;
assign ae_output_5b[4] = 5'b10010;
assign ae_output_5b[5] = 5'b10;
assign ae_output_5b[6] = 5'b0;
assign ae_output_5b[7] = 5'b11010;
assign ae_output_5b[8] = 5'b10101;
assign ae_output_5b[9] = 5'b10010;
assign ae_output_5b[10] = 5'b0;
assign ae_output_5b[11] = 5'b1;
assign ae_output_5b[12] = 5'b1;
assign ae_output_5b[13] = 5'b0;
assign ae_output_5b[14] = 5'b11111;
assign ae_output_5b[15] = 5'b11110;
assign ae_output_5b[16] = 5'b11111;
assign ae_output_5b[17] = 5'b1111;
assign ae_output_5b[18] = 5'b1;
assign ae_output_5b[19] = 5'b1;
assign ae_output_5b[20] = 5'b10;
assign ae_output_5b[21] = 5'b11;
assign ae_output_5b[22] = 5'b10101;
assign ae_output_5b[23] = 5'b10;
assign ae_output_5b[24] = 5'b11110;
assign ae_output_5b[25] = 5'b11110;
assign ae_output_5b[26] = 5'b10000;
assign ae_output_5b[27] = 5'b0;
assign ae_output_5b[28] = 5'b11101;
assign ae_output_5b[29] = 5'b10001;
// 7-bit output from original PCA weights (from Panpan)

assign pca_output_orig_7b[0] = 7'b1111111;
assign pca_output_orig_7b[1] = 7'b1111111;
assign pca_output_orig_7b[2] = 7'b0;
assign pca_output_orig_7b[3] = 7'b1111111;
assign pca_output_orig_7b[4] = 7'b0;
assign pca_output_orig_7b[5] = 7'b1111110;
assign pca_output_orig_7b[6] = 7'b1111111;
assign pca_output_orig_7b[7] = 7'b0;
assign pca_output_orig_7b[8] = 7'b0;
assign pca_output_orig_7b[9] = 7'b1111111;
assign pca_output_orig_7b[10] = 7'b1111111;
assign pca_output_orig_7b[11] = 7'b1111111;
assign pca_output_orig_7b[12] = 7'b1;
assign pca_output_orig_7b[13] = 7'b1;
assign pca_output_orig_7b[14] = 7'b1111011;
assign pca_output_orig_7b[15] = 7'b0;
assign pca_output_orig_7b[16] = 7'b1111110;
assign pca_output_orig_7b[17] = 7'b11;
assign pca_output_orig_7b[18] = 7'b1111101;
assign pca_output_orig_7b[19] = 7'b0;
assign pca_output_orig_7b[20] = 7'b1111101;
assign pca_output_orig_7b[21] = 7'b1111111;
assign pca_output_orig_7b[22] = 7'b1111110;
assign pca_output_orig_7b[23] = 7'b0;
assign pca_output_orig_7b[24] = 7'b1111111;
assign pca_output_orig_7b[25] = 7'b1111111;
assign pca_output_orig_7b[26] = 7'b1111111;
assign pca_output_orig_7b[27] = 7'b100;
assign pca_output_orig_7b[28] = 7'b1111100;
assign pca_output_orig_7b[29] = 7'b1111110;


